magic
tech sky130A
magscale 1 2
timestamp 1662591347
<< pwell >>
rect -1312 -1613 1312 1613
<< nmoslvt >>
rect -1116 865 -716 1465
rect -658 865 -258 1465
rect -200 865 200 1465
rect 258 865 658 1465
rect 716 865 1116 1465
rect -1116 109 -716 709
rect -658 109 -258 709
rect -200 109 200 709
rect 258 109 658 709
rect 716 109 1116 709
rect -1116 -647 -716 -47
rect -658 -647 -258 -47
rect -200 -647 200 -47
rect 258 -647 658 -47
rect 716 -647 1116 -47
rect -1116 -1403 -716 -803
rect -658 -1403 -258 -803
rect -200 -1403 200 -803
rect 258 -1403 658 -803
rect 716 -1403 1116 -803
<< ndiff >>
rect -1174 1453 -1116 1465
rect -1174 877 -1162 1453
rect -1128 877 -1116 1453
rect -1174 865 -1116 877
rect -716 1453 -658 1465
rect -716 877 -704 1453
rect -670 877 -658 1453
rect -716 865 -658 877
rect -258 1453 -200 1465
rect -258 877 -246 1453
rect -212 877 -200 1453
rect -258 865 -200 877
rect 200 1453 258 1465
rect 200 877 212 1453
rect 246 877 258 1453
rect 200 865 258 877
rect 658 1453 716 1465
rect 658 877 670 1453
rect 704 877 716 1453
rect 658 865 716 877
rect 1116 1453 1174 1465
rect 1116 877 1128 1453
rect 1162 877 1174 1453
rect 1116 865 1174 877
rect -1174 697 -1116 709
rect -1174 121 -1162 697
rect -1128 121 -1116 697
rect -1174 109 -1116 121
rect -716 697 -658 709
rect -716 121 -704 697
rect -670 121 -658 697
rect -716 109 -658 121
rect -258 697 -200 709
rect -258 121 -246 697
rect -212 121 -200 697
rect -258 109 -200 121
rect 200 697 258 709
rect 200 121 212 697
rect 246 121 258 697
rect 200 109 258 121
rect 658 697 716 709
rect 658 121 670 697
rect 704 121 716 697
rect 658 109 716 121
rect 1116 697 1174 709
rect 1116 121 1128 697
rect 1162 121 1174 697
rect 1116 109 1174 121
rect -1174 -59 -1116 -47
rect -1174 -635 -1162 -59
rect -1128 -635 -1116 -59
rect -1174 -647 -1116 -635
rect -716 -59 -658 -47
rect -716 -635 -704 -59
rect -670 -635 -658 -59
rect -716 -647 -658 -635
rect -258 -59 -200 -47
rect -258 -635 -246 -59
rect -212 -635 -200 -59
rect -258 -647 -200 -635
rect 200 -59 258 -47
rect 200 -635 212 -59
rect 246 -635 258 -59
rect 200 -647 258 -635
rect 658 -59 716 -47
rect 658 -635 670 -59
rect 704 -635 716 -59
rect 658 -647 716 -635
rect 1116 -59 1174 -47
rect 1116 -635 1128 -59
rect 1162 -635 1174 -59
rect 1116 -647 1174 -635
rect -1174 -815 -1116 -803
rect -1174 -1391 -1162 -815
rect -1128 -1391 -1116 -815
rect -1174 -1403 -1116 -1391
rect -716 -815 -658 -803
rect -716 -1391 -704 -815
rect -670 -1391 -658 -815
rect -716 -1403 -658 -1391
rect -258 -815 -200 -803
rect -258 -1391 -246 -815
rect -212 -1391 -200 -815
rect -258 -1403 -200 -1391
rect 200 -815 258 -803
rect 200 -1391 212 -815
rect 246 -1391 258 -815
rect 200 -1403 258 -1391
rect 658 -815 716 -803
rect 658 -1391 670 -815
rect 704 -1391 716 -815
rect 658 -1403 716 -1391
rect 1116 -815 1174 -803
rect 1116 -1391 1128 -815
rect 1162 -1391 1174 -815
rect 1116 -1403 1174 -1391
<< ndiffc >>
rect -1162 877 -1128 1453
rect -704 877 -670 1453
rect -246 877 -212 1453
rect 212 877 246 1453
rect 670 877 704 1453
rect 1128 877 1162 1453
rect -1162 121 -1128 697
rect -704 121 -670 697
rect -246 121 -212 697
rect 212 121 246 697
rect 670 121 704 697
rect 1128 121 1162 697
rect -1162 -635 -1128 -59
rect -704 -635 -670 -59
rect -246 -635 -212 -59
rect 212 -635 246 -59
rect 670 -635 704 -59
rect 1128 -635 1162 -59
rect -1162 -1391 -1128 -815
rect -704 -1391 -670 -815
rect -246 -1391 -212 -815
rect 212 -1391 246 -815
rect 670 -1391 704 -815
rect 1128 -1391 1162 -815
<< psubdiff >>
rect -1276 1543 -1180 1577
rect 1180 1543 1276 1577
rect -1276 -1543 -1242 1543
rect 1242 -1543 1276 1543
rect -1276 -1577 -1180 -1543
rect 1180 -1577 1276 -1543
<< psubdiffcont >>
rect -1180 1543 1180 1577
rect -1180 -1577 1180 -1543
<< poly >>
rect -1116 1465 -716 1491
rect -658 1465 -258 1491
rect -200 1465 200 1491
rect 258 1465 658 1491
rect 716 1465 1116 1491
rect -1116 827 -716 865
rect -1116 793 -1100 827
rect -732 793 -716 827
rect -1116 777 -716 793
rect -658 827 -258 865
rect -658 793 -642 827
rect -274 793 -258 827
rect -658 777 -258 793
rect -200 827 200 865
rect -200 793 -184 827
rect 184 793 200 827
rect -200 777 200 793
rect 258 827 658 865
rect 258 793 274 827
rect 642 793 658 827
rect 258 777 658 793
rect 716 827 1116 865
rect 716 793 732 827
rect 1100 793 1116 827
rect 716 777 1116 793
rect -1116 709 -716 735
rect -658 709 -258 735
rect -200 709 200 735
rect 258 709 658 735
rect 716 709 1116 735
rect -1116 71 -716 109
rect -1116 37 -1100 71
rect -732 37 -716 71
rect -1116 21 -716 37
rect -658 71 -258 109
rect -658 37 -642 71
rect -274 37 -258 71
rect -658 21 -258 37
rect -200 71 200 109
rect -200 37 -184 71
rect 184 37 200 71
rect -200 21 200 37
rect 258 71 658 109
rect 258 37 274 71
rect 642 37 658 71
rect 258 21 658 37
rect 716 71 1116 109
rect 716 37 732 71
rect 1100 37 1116 71
rect 716 21 1116 37
rect -1116 -47 -716 -21
rect -658 -47 -258 -21
rect -200 -47 200 -21
rect 258 -47 658 -21
rect 716 -47 1116 -21
rect -1116 -685 -716 -647
rect -1116 -719 -1100 -685
rect -732 -719 -716 -685
rect -1116 -735 -716 -719
rect -658 -685 -258 -647
rect -658 -719 -642 -685
rect -274 -719 -258 -685
rect -658 -735 -258 -719
rect -200 -685 200 -647
rect -200 -719 -184 -685
rect 184 -719 200 -685
rect -200 -735 200 -719
rect 258 -685 658 -647
rect 258 -719 274 -685
rect 642 -719 658 -685
rect 258 -735 658 -719
rect 716 -685 1116 -647
rect 716 -719 732 -685
rect 1100 -719 1116 -685
rect 716 -735 1116 -719
rect -1116 -803 -716 -777
rect -658 -803 -258 -777
rect -200 -803 200 -777
rect 258 -803 658 -777
rect 716 -803 1116 -777
rect -1116 -1441 -716 -1403
rect -1116 -1475 -1100 -1441
rect -732 -1475 -716 -1441
rect -1116 -1491 -716 -1475
rect -658 -1441 -258 -1403
rect -658 -1475 -642 -1441
rect -274 -1475 -258 -1441
rect -658 -1491 -258 -1475
rect -200 -1441 200 -1403
rect -200 -1475 -184 -1441
rect 184 -1475 200 -1441
rect -200 -1491 200 -1475
rect 258 -1441 658 -1403
rect 258 -1475 274 -1441
rect 642 -1475 658 -1441
rect 258 -1491 658 -1475
rect 716 -1441 1116 -1403
rect 716 -1475 732 -1441
rect 1100 -1475 1116 -1441
rect 716 -1491 1116 -1475
<< polycont >>
rect -1100 793 -732 827
rect -642 793 -274 827
rect -184 793 184 827
rect 274 793 642 827
rect 732 793 1100 827
rect -1100 37 -732 71
rect -642 37 -274 71
rect -184 37 184 71
rect 274 37 642 71
rect 732 37 1100 71
rect -1100 -719 -732 -685
rect -642 -719 -274 -685
rect -184 -719 184 -685
rect 274 -719 642 -685
rect 732 -719 1100 -685
rect -1100 -1475 -732 -1441
rect -642 -1475 -274 -1441
rect -184 -1475 184 -1441
rect 274 -1475 642 -1441
rect 732 -1475 1100 -1441
<< locali >>
rect -1276 1543 -1180 1577
rect 1180 1543 1276 1577
rect -1276 -1543 -1242 1543
rect -1162 1453 -1128 1469
rect -1162 861 -1128 877
rect -704 1453 -670 1469
rect -704 861 -670 877
rect -246 1453 -212 1469
rect -246 861 -212 877
rect 212 1453 246 1469
rect 212 861 246 877
rect 670 1453 704 1469
rect 670 861 704 877
rect 1128 1453 1162 1469
rect 1128 861 1162 877
rect -1116 793 -1100 827
rect -732 793 -716 827
rect -658 793 -642 827
rect -274 793 -258 827
rect -200 793 -184 827
rect 184 793 200 827
rect 258 793 274 827
rect 642 793 658 827
rect 716 793 732 827
rect 1100 793 1116 827
rect -1162 697 -1128 713
rect -1162 105 -1128 121
rect -704 697 -670 713
rect -704 105 -670 121
rect -246 697 -212 713
rect -246 105 -212 121
rect 212 697 246 713
rect 212 105 246 121
rect 670 697 704 713
rect 670 105 704 121
rect 1128 697 1162 713
rect 1128 105 1162 121
rect -1116 37 -1100 71
rect -732 37 -716 71
rect -658 37 -642 71
rect -274 37 -258 71
rect -200 37 -184 71
rect 184 37 200 71
rect 258 37 274 71
rect 642 37 658 71
rect 716 37 732 71
rect 1100 37 1116 71
rect -1162 -59 -1128 -43
rect -1162 -651 -1128 -635
rect -704 -59 -670 -43
rect -704 -651 -670 -635
rect -246 -59 -212 -43
rect -246 -651 -212 -635
rect 212 -59 246 -43
rect 212 -651 246 -635
rect 670 -59 704 -43
rect 670 -651 704 -635
rect 1128 -59 1162 -43
rect 1128 -651 1162 -635
rect -1116 -719 -1100 -685
rect -732 -719 -716 -685
rect -658 -719 -642 -685
rect -274 -719 -258 -685
rect -200 -719 -184 -685
rect 184 -719 200 -685
rect 258 -719 274 -685
rect 642 -719 658 -685
rect 716 -719 732 -685
rect 1100 -719 1116 -685
rect -1162 -815 -1128 -799
rect -1162 -1407 -1128 -1391
rect -704 -815 -670 -799
rect -704 -1407 -670 -1391
rect -246 -815 -212 -799
rect -246 -1407 -212 -1391
rect 212 -815 246 -799
rect 212 -1407 246 -1391
rect 670 -815 704 -799
rect 670 -1407 704 -1391
rect 1128 -815 1162 -799
rect 1128 -1407 1162 -1391
rect -1116 -1475 -1100 -1441
rect -732 -1475 -716 -1441
rect -658 -1475 -642 -1441
rect -274 -1475 -258 -1441
rect -200 -1475 -184 -1441
rect 184 -1475 200 -1441
rect 258 -1475 274 -1441
rect 642 -1475 658 -1441
rect 716 -1475 732 -1441
rect 1100 -1475 1116 -1441
rect 1242 -1543 1276 1543
rect -1276 -1577 -1180 -1543
rect 1180 -1577 1276 -1543
<< viali >>
rect -1162 877 -1128 1453
rect -704 877 -670 1453
rect -246 877 -212 1453
rect 212 877 246 1453
rect 670 877 704 1453
rect 1128 877 1162 1453
rect -1100 793 -732 827
rect -642 793 -274 827
rect -184 793 184 827
rect 274 793 642 827
rect 732 793 1100 827
rect -1162 121 -1128 697
rect -704 121 -670 697
rect -246 121 -212 697
rect 212 121 246 697
rect 670 121 704 697
rect 1128 121 1162 697
rect -1100 37 -732 71
rect -642 37 -274 71
rect -184 37 184 71
rect 274 37 642 71
rect 732 37 1100 71
rect -1162 -635 -1128 -59
rect -704 -635 -670 -59
rect -246 -635 -212 -59
rect 212 -635 246 -59
rect 670 -635 704 -59
rect 1128 -635 1162 -59
rect -1100 -719 -732 -685
rect -642 -719 -274 -685
rect -184 -719 184 -685
rect 274 -719 642 -685
rect 732 -719 1100 -685
rect -1162 -1391 -1128 -815
rect -704 -1391 -670 -815
rect -246 -1391 -212 -815
rect 212 -1391 246 -815
rect 670 -1391 704 -815
rect 1128 -1391 1162 -815
rect -1100 -1475 -732 -1441
rect -642 -1475 -274 -1441
rect -184 -1475 184 -1441
rect 274 -1475 642 -1441
rect 732 -1475 1100 -1441
<< metal1 >>
rect -1168 1453 -1122 1465
rect -1168 877 -1162 1453
rect -1128 877 -1122 1453
rect -1168 865 -1122 877
rect -710 1453 -664 1465
rect -710 877 -704 1453
rect -670 877 -664 1453
rect -710 865 -664 877
rect -252 1453 -206 1465
rect -252 877 -246 1453
rect -212 877 -206 1453
rect -252 865 -206 877
rect 206 1453 252 1465
rect 206 877 212 1453
rect 246 877 252 1453
rect 206 865 252 877
rect 664 1453 710 1465
rect 664 877 670 1453
rect 704 877 710 1453
rect 664 865 710 877
rect 1122 1453 1168 1465
rect 1122 877 1128 1453
rect 1162 877 1168 1453
rect 1122 865 1168 877
rect -1112 827 -720 833
rect -1112 793 -1100 827
rect -732 793 -720 827
rect -1112 787 -720 793
rect -654 827 -262 833
rect -654 793 -642 827
rect -274 793 -262 827
rect -654 787 -262 793
rect -196 827 196 833
rect -196 793 -184 827
rect 184 793 196 827
rect -196 787 196 793
rect 262 827 654 833
rect 262 793 274 827
rect 642 793 654 827
rect 262 787 654 793
rect 720 827 1112 833
rect 720 793 732 827
rect 1100 793 1112 827
rect 720 787 1112 793
rect -1168 697 -1122 709
rect -1168 121 -1162 697
rect -1128 121 -1122 697
rect -1168 109 -1122 121
rect -710 697 -664 709
rect -710 121 -704 697
rect -670 121 -664 697
rect -710 109 -664 121
rect -252 697 -206 709
rect -252 121 -246 697
rect -212 121 -206 697
rect -252 109 -206 121
rect 206 697 252 709
rect 206 121 212 697
rect 246 121 252 697
rect 206 109 252 121
rect 664 697 710 709
rect 664 121 670 697
rect 704 121 710 697
rect 664 109 710 121
rect 1122 697 1168 709
rect 1122 121 1128 697
rect 1162 121 1168 697
rect 1122 109 1168 121
rect -1112 71 -720 77
rect -1112 37 -1100 71
rect -732 37 -720 71
rect -1112 31 -720 37
rect -654 71 -262 77
rect -654 37 -642 71
rect -274 37 -262 71
rect -654 31 -262 37
rect -196 71 196 77
rect -196 37 -184 71
rect 184 37 196 71
rect -196 31 196 37
rect 262 71 654 77
rect 262 37 274 71
rect 642 37 654 71
rect 262 31 654 37
rect 720 71 1112 77
rect 720 37 732 71
rect 1100 37 1112 71
rect 720 31 1112 37
rect -1168 -59 -1122 -47
rect -1168 -635 -1162 -59
rect -1128 -635 -1122 -59
rect -1168 -647 -1122 -635
rect -710 -59 -664 -47
rect -710 -635 -704 -59
rect -670 -635 -664 -59
rect -710 -647 -664 -635
rect -252 -59 -206 -47
rect -252 -635 -246 -59
rect -212 -635 -206 -59
rect -252 -647 -206 -635
rect 206 -59 252 -47
rect 206 -635 212 -59
rect 246 -635 252 -59
rect 206 -647 252 -635
rect 664 -59 710 -47
rect 664 -635 670 -59
rect 704 -635 710 -59
rect 664 -647 710 -635
rect 1122 -59 1168 -47
rect 1122 -635 1128 -59
rect 1162 -635 1168 -59
rect 1122 -647 1168 -635
rect -1112 -685 -720 -679
rect -1112 -719 -1100 -685
rect -732 -719 -720 -685
rect -1112 -725 -720 -719
rect -654 -685 -262 -679
rect -654 -719 -642 -685
rect -274 -719 -262 -685
rect -654 -725 -262 -719
rect -196 -685 196 -679
rect -196 -719 -184 -685
rect 184 -719 196 -685
rect -196 -725 196 -719
rect 262 -685 654 -679
rect 262 -719 274 -685
rect 642 -719 654 -685
rect 262 -725 654 -719
rect 720 -685 1112 -679
rect 720 -719 732 -685
rect 1100 -719 1112 -685
rect 720 -725 1112 -719
rect -1168 -815 -1122 -803
rect -1168 -1391 -1162 -815
rect -1128 -1391 -1122 -815
rect -1168 -1403 -1122 -1391
rect -710 -815 -664 -803
rect -710 -1391 -704 -815
rect -670 -1391 -664 -815
rect -710 -1403 -664 -1391
rect -252 -815 -206 -803
rect -252 -1391 -246 -815
rect -212 -1391 -206 -815
rect -252 -1403 -206 -1391
rect 206 -815 252 -803
rect 206 -1391 212 -815
rect 246 -1391 252 -815
rect 206 -1403 252 -1391
rect 664 -815 710 -803
rect 664 -1391 670 -815
rect 704 -1391 710 -815
rect 664 -1403 710 -1391
rect 1122 -815 1168 -803
rect 1122 -1391 1128 -815
rect 1162 -1391 1168 -815
rect 1122 -1403 1168 -1391
rect -1112 -1441 -720 -1435
rect -1112 -1475 -1100 -1441
rect -732 -1475 -720 -1441
rect -1112 -1481 -720 -1475
rect -654 -1441 -262 -1435
rect -654 -1475 -642 -1441
rect -274 -1475 -262 -1441
rect -654 -1481 -262 -1475
rect -196 -1441 196 -1435
rect -196 -1475 -184 -1441
rect 184 -1475 196 -1441
rect -196 -1481 196 -1475
rect 262 -1441 654 -1435
rect 262 -1475 274 -1441
rect 642 -1475 654 -1441
rect 262 -1481 654 -1475
rect 720 -1441 1112 -1435
rect 720 -1475 732 -1441
rect 1100 -1475 1112 -1441
rect 720 -1481 1112 -1475
<< properties >>
string FIXED_BBOX -1259 -1560 1259 1560
string gencell sky130_fd_pr__nfet_01v8_lvt
string library sky130
string parameters w 3 l 2 m 4 nf 5 diffcov 100 polycov 100 guard 1 glc 0 grc 0 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 0 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
