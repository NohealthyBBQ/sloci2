magic
tech sky130A
magscale 1 2
timestamp 1662671450
<< nwell >>
rect -296 -6205 296 6205
<< pmoslvt >>
rect -100 5786 100 5986
rect -100 5350 100 5550
rect -100 4914 100 5114
rect -100 4478 100 4678
rect -100 4042 100 4242
rect -100 3606 100 3806
rect -100 3170 100 3370
rect -100 2734 100 2934
rect -100 2298 100 2498
rect -100 1862 100 2062
rect -100 1426 100 1626
rect -100 990 100 1190
rect -100 554 100 754
rect -100 118 100 318
rect -100 -318 100 -118
rect -100 -754 100 -554
rect -100 -1190 100 -990
rect -100 -1626 100 -1426
rect -100 -2062 100 -1862
rect -100 -2498 100 -2298
rect -100 -2934 100 -2734
rect -100 -3370 100 -3170
rect -100 -3806 100 -3606
rect -100 -4242 100 -4042
rect -100 -4678 100 -4478
rect -100 -5114 100 -4914
rect -100 -5550 100 -5350
rect -100 -5986 100 -5786
<< pdiff >>
rect -158 5974 -100 5986
rect -158 5798 -146 5974
rect -112 5798 -100 5974
rect -158 5786 -100 5798
rect 100 5974 158 5986
rect 100 5798 112 5974
rect 146 5798 158 5974
rect 100 5786 158 5798
rect -158 5538 -100 5550
rect -158 5362 -146 5538
rect -112 5362 -100 5538
rect -158 5350 -100 5362
rect 100 5538 158 5550
rect 100 5362 112 5538
rect 146 5362 158 5538
rect 100 5350 158 5362
rect -158 5102 -100 5114
rect -158 4926 -146 5102
rect -112 4926 -100 5102
rect -158 4914 -100 4926
rect 100 5102 158 5114
rect 100 4926 112 5102
rect 146 4926 158 5102
rect 100 4914 158 4926
rect -158 4666 -100 4678
rect -158 4490 -146 4666
rect -112 4490 -100 4666
rect -158 4478 -100 4490
rect 100 4666 158 4678
rect 100 4490 112 4666
rect 146 4490 158 4666
rect 100 4478 158 4490
rect -158 4230 -100 4242
rect -158 4054 -146 4230
rect -112 4054 -100 4230
rect -158 4042 -100 4054
rect 100 4230 158 4242
rect 100 4054 112 4230
rect 146 4054 158 4230
rect 100 4042 158 4054
rect -158 3794 -100 3806
rect -158 3618 -146 3794
rect -112 3618 -100 3794
rect -158 3606 -100 3618
rect 100 3794 158 3806
rect 100 3618 112 3794
rect 146 3618 158 3794
rect 100 3606 158 3618
rect -158 3358 -100 3370
rect -158 3182 -146 3358
rect -112 3182 -100 3358
rect -158 3170 -100 3182
rect 100 3358 158 3370
rect 100 3182 112 3358
rect 146 3182 158 3358
rect 100 3170 158 3182
rect -158 2922 -100 2934
rect -158 2746 -146 2922
rect -112 2746 -100 2922
rect -158 2734 -100 2746
rect 100 2922 158 2934
rect 100 2746 112 2922
rect 146 2746 158 2922
rect 100 2734 158 2746
rect -158 2486 -100 2498
rect -158 2310 -146 2486
rect -112 2310 -100 2486
rect -158 2298 -100 2310
rect 100 2486 158 2498
rect 100 2310 112 2486
rect 146 2310 158 2486
rect 100 2298 158 2310
rect -158 2050 -100 2062
rect -158 1874 -146 2050
rect -112 1874 -100 2050
rect -158 1862 -100 1874
rect 100 2050 158 2062
rect 100 1874 112 2050
rect 146 1874 158 2050
rect 100 1862 158 1874
rect -158 1614 -100 1626
rect -158 1438 -146 1614
rect -112 1438 -100 1614
rect -158 1426 -100 1438
rect 100 1614 158 1626
rect 100 1438 112 1614
rect 146 1438 158 1614
rect 100 1426 158 1438
rect -158 1178 -100 1190
rect -158 1002 -146 1178
rect -112 1002 -100 1178
rect -158 990 -100 1002
rect 100 1178 158 1190
rect 100 1002 112 1178
rect 146 1002 158 1178
rect 100 990 158 1002
rect -158 742 -100 754
rect -158 566 -146 742
rect -112 566 -100 742
rect -158 554 -100 566
rect 100 742 158 754
rect 100 566 112 742
rect 146 566 158 742
rect 100 554 158 566
rect -158 306 -100 318
rect -158 130 -146 306
rect -112 130 -100 306
rect -158 118 -100 130
rect 100 306 158 318
rect 100 130 112 306
rect 146 130 158 306
rect 100 118 158 130
rect -158 -130 -100 -118
rect -158 -306 -146 -130
rect -112 -306 -100 -130
rect -158 -318 -100 -306
rect 100 -130 158 -118
rect 100 -306 112 -130
rect 146 -306 158 -130
rect 100 -318 158 -306
rect -158 -566 -100 -554
rect -158 -742 -146 -566
rect -112 -742 -100 -566
rect -158 -754 -100 -742
rect 100 -566 158 -554
rect 100 -742 112 -566
rect 146 -742 158 -566
rect 100 -754 158 -742
rect -158 -1002 -100 -990
rect -158 -1178 -146 -1002
rect -112 -1178 -100 -1002
rect -158 -1190 -100 -1178
rect 100 -1002 158 -990
rect 100 -1178 112 -1002
rect 146 -1178 158 -1002
rect 100 -1190 158 -1178
rect -158 -1438 -100 -1426
rect -158 -1614 -146 -1438
rect -112 -1614 -100 -1438
rect -158 -1626 -100 -1614
rect 100 -1438 158 -1426
rect 100 -1614 112 -1438
rect 146 -1614 158 -1438
rect 100 -1626 158 -1614
rect -158 -1874 -100 -1862
rect -158 -2050 -146 -1874
rect -112 -2050 -100 -1874
rect -158 -2062 -100 -2050
rect 100 -1874 158 -1862
rect 100 -2050 112 -1874
rect 146 -2050 158 -1874
rect 100 -2062 158 -2050
rect -158 -2310 -100 -2298
rect -158 -2486 -146 -2310
rect -112 -2486 -100 -2310
rect -158 -2498 -100 -2486
rect 100 -2310 158 -2298
rect 100 -2486 112 -2310
rect 146 -2486 158 -2310
rect 100 -2498 158 -2486
rect -158 -2746 -100 -2734
rect -158 -2922 -146 -2746
rect -112 -2922 -100 -2746
rect -158 -2934 -100 -2922
rect 100 -2746 158 -2734
rect 100 -2922 112 -2746
rect 146 -2922 158 -2746
rect 100 -2934 158 -2922
rect -158 -3182 -100 -3170
rect -158 -3358 -146 -3182
rect -112 -3358 -100 -3182
rect -158 -3370 -100 -3358
rect 100 -3182 158 -3170
rect 100 -3358 112 -3182
rect 146 -3358 158 -3182
rect 100 -3370 158 -3358
rect -158 -3618 -100 -3606
rect -158 -3794 -146 -3618
rect -112 -3794 -100 -3618
rect -158 -3806 -100 -3794
rect 100 -3618 158 -3606
rect 100 -3794 112 -3618
rect 146 -3794 158 -3618
rect 100 -3806 158 -3794
rect -158 -4054 -100 -4042
rect -158 -4230 -146 -4054
rect -112 -4230 -100 -4054
rect -158 -4242 -100 -4230
rect 100 -4054 158 -4042
rect 100 -4230 112 -4054
rect 146 -4230 158 -4054
rect 100 -4242 158 -4230
rect -158 -4490 -100 -4478
rect -158 -4666 -146 -4490
rect -112 -4666 -100 -4490
rect -158 -4678 -100 -4666
rect 100 -4490 158 -4478
rect 100 -4666 112 -4490
rect 146 -4666 158 -4490
rect 100 -4678 158 -4666
rect -158 -4926 -100 -4914
rect -158 -5102 -146 -4926
rect -112 -5102 -100 -4926
rect -158 -5114 -100 -5102
rect 100 -4926 158 -4914
rect 100 -5102 112 -4926
rect 146 -5102 158 -4926
rect 100 -5114 158 -5102
rect -158 -5362 -100 -5350
rect -158 -5538 -146 -5362
rect -112 -5538 -100 -5362
rect -158 -5550 -100 -5538
rect 100 -5362 158 -5350
rect 100 -5538 112 -5362
rect 146 -5538 158 -5362
rect 100 -5550 158 -5538
rect -158 -5798 -100 -5786
rect -158 -5974 -146 -5798
rect -112 -5974 -100 -5798
rect -158 -5986 -100 -5974
rect 100 -5798 158 -5786
rect 100 -5974 112 -5798
rect 146 -5974 158 -5798
rect 100 -5986 158 -5974
<< pdiffc >>
rect -146 5798 -112 5974
rect 112 5798 146 5974
rect -146 5362 -112 5538
rect 112 5362 146 5538
rect -146 4926 -112 5102
rect 112 4926 146 5102
rect -146 4490 -112 4666
rect 112 4490 146 4666
rect -146 4054 -112 4230
rect 112 4054 146 4230
rect -146 3618 -112 3794
rect 112 3618 146 3794
rect -146 3182 -112 3358
rect 112 3182 146 3358
rect -146 2746 -112 2922
rect 112 2746 146 2922
rect -146 2310 -112 2486
rect 112 2310 146 2486
rect -146 1874 -112 2050
rect 112 1874 146 2050
rect -146 1438 -112 1614
rect 112 1438 146 1614
rect -146 1002 -112 1178
rect 112 1002 146 1178
rect -146 566 -112 742
rect 112 566 146 742
rect -146 130 -112 306
rect 112 130 146 306
rect -146 -306 -112 -130
rect 112 -306 146 -130
rect -146 -742 -112 -566
rect 112 -742 146 -566
rect -146 -1178 -112 -1002
rect 112 -1178 146 -1002
rect -146 -1614 -112 -1438
rect 112 -1614 146 -1438
rect -146 -2050 -112 -1874
rect 112 -2050 146 -1874
rect -146 -2486 -112 -2310
rect 112 -2486 146 -2310
rect -146 -2922 -112 -2746
rect 112 -2922 146 -2746
rect -146 -3358 -112 -3182
rect 112 -3358 146 -3182
rect -146 -3794 -112 -3618
rect 112 -3794 146 -3618
rect -146 -4230 -112 -4054
rect 112 -4230 146 -4054
rect -146 -4666 -112 -4490
rect 112 -4666 146 -4490
rect -146 -5102 -112 -4926
rect 112 -5102 146 -4926
rect -146 -5538 -112 -5362
rect 112 -5538 146 -5362
rect -146 -5974 -112 -5798
rect 112 -5974 146 -5798
<< nsubdiff >>
rect -260 6135 -164 6169
rect 164 6135 260 6169
rect -260 6073 -226 6135
rect 226 6073 260 6135
rect -260 -6135 -226 -6073
rect 226 -6135 260 -6073
rect -260 -6169 -164 -6135
rect 164 -6169 260 -6135
<< nsubdiffcont >>
rect -164 6135 164 6169
rect -260 -6073 -226 6073
rect 226 -6073 260 6073
rect -164 -6169 164 -6135
<< poly >>
rect -100 6067 100 6083
rect -100 6033 -84 6067
rect 84 6033 100 6067
rect -100 5986 100 6033
rect -100 5739 100 5786
rect -100 5705 -84 5739
rect 84 5705 100 5739
rect -100 5689 100 5705
rect -100 5631 100 5647
rect -100 5597 -84 5631
rect 84 5597 100 5631
rect -100 5550 100 5597
rect -100 5303 100 5350
rect -100 5269 -84 5303
rect 84 5269 100 5303
rect -100 5253 100 5269
rect -100 5195 100 5211
rect -100 5161 -84 5195
rect 84 5161 100 5195
rect -100 5114 100 5161
rect -100 4867 100 4914
rect -100 4833 -84 4867
rect 84 4833 100 4867
rect -100 4817 100 4833
rect -100 4759 100 4775
rect -100 4725 -84 4759
rect 84 4725 100 4759
rect -100 4678 100 4725
rect -100 4431 100 4478
rect -100 4397 -84 4431
rect 84 4397 100 4431
rect -100 4381 100 4397
rect -100 4323 100 4339
rect -100 4289 -84 4323
rect 84 4289 100 4323
rect -100 4242 100 4289
rect -100 3995 100 4042
rect -100 3961 -84 3995
rect 84 3961 100 3995
rect -100 3945 100 3961
rect -100 3887 100 3903
rect -100 3853 -84 3887
rect 84 3853 100 3887
rect -100 3806 100 3853
rect -100 3559 100 3606
rect -100 3525 -84 3559
rect 84 3525 100 3559
rect -100 3509 100 3525
rect -100 3451 100 3467
rect -100 3417 -84 3451
rect 84 3417 100 3451
rect -100 3370 100 3417
rect -100 3123 100 3170
rect -100 3089 -84 3123
rect 84 3089 100 3123
rect -100 3073 100 3089
rect -100 3015 100 3031
rect -100 2981 -84 3015
rect 84 2981 100 3015
rect -100 2934 100 2981
rect -100 2687 100 2734
rect -100 2653 -84 2687
rect 84 2653 100 2687
rect -100 2637 100 2653
rect -100 2579 100 2595
rect -100 2545 -84 2579
rect 84 2545 100 2579
rect -100 2498 100 2545
rect -100 2251 100 2298
rect -100 2217 -84 2251
rect 84 2217 100 2251
rect -100 2201 100 2217
rect -100 2143 100 2159
rect -100 2109 -84 2143
rect 84 2109 100 2143
rect -100 2062 100 2109
rect -100 1815 100 1862
rect -100 1781 -84 1815
rect 84 1781 100 1815
rect -100 1765 100 1781
rect -100 1707 100 1723
rect -100 1673 -84 1707
rect 84 1673 100 1707
rect -100 1626 100 1673
rect -100 1379 100 1426
rect -100 1345 -84 1379
rect 84 1345 100 1379
rect -100 1329 100 1345
rect -100 1271 100 1287
rect -100 1237 -84 1271
rect 84 1237 100 1271
rect -100 1190 100 1237
rect -100 943 100 990
rect -100 909 -84 943
rect 84 909 100 943
rect -100 893 100 909
rect -100 835 100 851
rect -100 801 -84 835
rect 84 801 100 835
rect -100 754 100 801
rect -100 507 100 554
rect -100 473 -84 507
rect 84 473 100 507
rect -100 457 100 473
rect -100 399 100 415
rect -100 365 -84 399
rect 84 365 100 399
rect -100 318 100 365
rect -100 71 100 118
rect -100 37 -84 71
rect 84 37 100 71
rect -100 21 100 37
rect -100 -37 100 -21
rect -100 -71 -84 -37
rect 84 -71 100 -37
rect -100 -118 100 -71
rect -100 -365 100 -318
rect -100 -399 -84 -365
rect 84 -399 100 -365
rect -100 -415 100 -399
rect -100 -473 100 -457
rect -100 -507 -84 -473
rect 84 -507 100 -473
rect -100 -554 100 -507
rect -100 -801 100 -754
rect -100 -835 -84 -801
rect 84 -835 100 -801
rect -100 -851 100 -835
rect -100 -909 100 -893
rect -100 -943 -84 -909
rect 84 -943 100 -909
rect -100 -990 100 -943
rect -100 -1237 100 -1190
rect -100 -1271 -84 -1237
rect 84 -1271 100 -1237
rect -100 -1287 100 -1271
rect -100 -1345 100 -1329
rect -100 -1379 -84 -1345
rect 84 -1379 100 -1345
rect -100 -1426 100 -1379
rect -100 -1673 100 -1626
rect -100 -1707 -84 -1673
rect 84 -1707 100 -1673
rect -100 -1723 100 -1707
rect -100 -1781 100 -1765
rect -100 -1815 -84 -1781
rect 84 -1815 100 -1781
rect -100 -1862 100 -1815
rect -100 -2109 100 -2062
rect -100 -2143 -84 -2109
rect 84 -2143 100 -2109
rect -100 -2159 100 -2143
rect -100 -2217 100 -2201
rect -100 -2251 -84 -2217
rect 84 -2251 100 -2217
rect -100 -2298 100 -2251
rect -100 -2545 100 -2498
rect -100 -2579 -84 -2545
rect 84 -2579 100 -2545
rect -100 -2595 100 -2579
rect -100 -2653 100 -2637
rect -100 -2687 -84 -2653
rect 84 -2687 100 -2653
rect -100 -2734 100 -2687
rect -100 -2981 100 -2934
rect -100 -3015 -84 -2981
rect 84 -3015 100 -2981
rect -100 -3031 100 -3015
rect -100 -3089 100 -3073
rect -100 -3123 -84 -3089
rect 84 -3123 100 -3089
rect -100 -3170 100 -3123
rect -100 -3417 100 -3370
rect -100 -3451 -84 -3417
rect 84 -3451 100 -3417
rect -100 -3467 100 -3451
rect -100 -3525 100 -3509
rect -100 -3559 -84 -3525
rect 84 -3559 100 -3525
rect -100 -3606 100 -3559
rect -100 -3853 100 -3806
rect -100 -3887 -84 -3853
rect 84 -3887 100 -3853
rect -100 -3903 100 -3887
rect -100 -3961 100 -3945
rect -100 -3995 -84 -3961
rect 84 -3995 100 -3961
rect -100 -4042 100 -3995
rect -100 -4289 100 -4242
rect -100 -4323 -84 -4289
rect 84 -4323 100 -4289
rect -100 -4339 100 -4323
rect -100 -4397 100 -4381
rect -100 -4431 -84 -4397
rect 84 -4431 100 -4397
rect -100 -4478 100 -4431
rect -100 -4725 100 -4678
rect -100 -4759 -84 -4725
rect 84 -4759 100 -4725
rect -100 -4775 100 -4759
rect -100 -4833 100 -4817
rect -100 -4867 -84 -4833
rect 84 -4867 100 -4833
rect -100 -4914 100 -4867
rect -100 -5161 100 -5114
rect -100 -5195 -84 -5161
rect 84 -5195 100 -5161
rect -100 -5211 100 -5195
rect -100 -5269 100 -5253
rect -100 -5303 -84 -5269
rect 84 -5303 100 -5269
rect -100 -5350 100 -5303
rect -100 -5597 100 -5550
rect -100 -5631 -84 -5597
rect 84 -5631 100 -5597
rect -100 -5647 100 -5631
rect -100 -5705 100 -5689
rect -100 -5739 -84 -5705
rect 84 -5739 100 -5705
rect -100 -5786 100 -5739
rect -100 -6033 100 -5986
rect -100 -6067 -84 -6033
rect 84 -6067 100 -6033
rect -100 -6083 100 -6067
<< polycont >>
rect -84 6033 84 6067
rect -84 5705 84 5739
rect -84 5597 84 5631
rect -84 5269 84 5303
rect -84 5161 84 5195
rect -84 4833 84 4867
rect -84 4725 84 4759
rect -84 4397 84 4431
rect -84 4289 84 4323
rect -84 3961 84 3995
rect -84 3853 84 3887
rect -84 3525 84 3559
rect -84 3417 84 3451
rect -84 3089 84 3123
rect -84 2981 84 3015
rect -84 2653 84 2687
rect -84 2545 84 2579
rect -84 2217 84 2251
rect -84 2109 84 2143
rect -84 1781 84 1815
rect -84 1673 84 1707
rect -84 1345 84 1379
rect -84 1237 84 1271
rect -84 909 84 943
rect -84 801 84 835
rect -84 473 84 507
rect -84 365 84 399
rect -84 37 84 71
rect -84 -71 84 -37
rect -84 -399 84 -365
rect -84 -507 84 -473
rect -84 -835 84 -801
rect -84 -943 84 -909
rect -84 -1271 84 -1237
rect -84 -1379 84 -1345
rect -84 -1707 84 -1673
rect -84 -1815 84 -1781
rect -84 -2143 84 -2109
rect -84 -2251 84 -2217
rect -84 -2579 84 -2545
rect -84 -2687 84 -2653
rect -84 -3015 84 -2981
rect -84 -3123 84 -3089
rect -84 -3451 84 -3417
rect -84 -3559 84 -3525
rect -84 -3887 84 -3853
rect -84 -3995 84 -3961
rect -84 -4323 84 -4289
rect -84 -4431 84 -4397
rect -84 -4759 84 -4725
rect -84 -4867 84 -4833
rect -84 -5195 84 -5161
rect -84 -5303 84 -5269
rect -84 -5631 84 -5597
rect -84 -5739 84 -5705
rect -84 -6067 84 -6033
<< locali >>
rect -260 6135 -164 6169
rect 164 6135 260 6169
rect -260 6073 -226 6135
rect 226 6073 260 6135
rect -100 6033 -84 6067
rect 84 6033 100 6067
rect -146 5974 -112 5990
rect -146 5782 -112 5798
rect 112 5974 146 5990
rect 112 5782 146 5798
rect -100 5705 -84 5739
rect 84 5705 100 5739
rect -100 5597 -84 5631
rect 84 5597 100 5631
rect -146 5538 -112 5554
rect -146 5346 -112 5362
rect 112 5538 146 5554
rect 112 5346 146 5362
rect -100 5269 -84 5303
rect 84 5269 100 5303
rect -100 5161 -84 5195
rect 84 5161 100 5195
rect -146 5102 -112 5118
rect -146 4910 -112 4926
rect 112 5102 146 5118
rect 112 4910 146 4926
rect -100 4833 -84 4867
rect 84 4833 100 4867
rect -100 4725 -84 4759
rect 84 4725 100 4759
rect -146 4666 -112 4682
rect -146 4474 -112 4490
rect 112 4666 146 4682
rect 112 4474 146 4490
rect -100 4397 -84 4431
rect 84 4397 100 4431
rect -100 4289 -84 4323
rect 84 4289 100 4323
rect -146 4230 -112 4246
rect -146 4038 -112 4054
rect 112 4230 146 4246
rect 112 4038 146 4054
rect -100 3961 -84 3995
rect 84 3961 100 3995
rect -100 3853 -84 3887
rect 84 3853 100 3887
rect -146 3794 -112 3810
rect -146 3602 -112 3618
rect 112 3794 146 3810
rect 112 3602 146 3618
rect -100 3525 -84 3559
rect 84 3525 100 3559
rect -100 3417 -84 3451
rect 84 3417 100 3451
rect -146 3358 -112 3374
rect -146 3166 -112 3182
rect 112 3358 146 3374
rect 112 3166 146 3182
rect -100 3089 -84 3123
rect 84 3089 100 3123
rect -100 2981 -84 3015
rect 84 2981 100 3015
rect -146 2922 -112 2938
rect -146 2730 -112 2746
rect 112 2922 146 2938
rect 112 2730 146 2746
rect -100 2653 -84 2687
rect 84 2653 100 2687
rect -100 2545 -84 2579
rect 84 2545 100 2579
rect -146 2486 -112 2502
rect -146 2294 -112 2310
rect 112 2486 146 2502
rect 112 2294 146 2310
rect -100 2217 -84 2251
rect 84 2217 100 2251
rect -100 2109 -84 2143
rect 84 2109 100 2143
rect -146 2050 -112 2066
rect -146 1858 -112 1874
rect 112 2050 146 2066
rect 112 1858 146 1874
rect -100 1781 -84 1815
rect 84 1781 100 1815
rect -100 1673 -84 1707
rect 84 1673 100 1707
rect -146 1614 -112 1630
rect -146 1422 -112 1438
rect 112 1614 146 1630
rect 112 1422 146 1438
rect -100 1345 -84 1379
rect 84 1345 100 1379
rect -100 1237 -84 1271
rect 84 1237 100 1271
rect -146 1178 -112 1194
rect -146 986 -112 1002
rect 112 1178 146 1194
rect 112 986 146 1002
rect -100 909 -84 943
rect 84 909 100 943
rect -100 801 -84 835
rect 84 801 100 835
rect -146 742 -112 758
rect -146 550 -112 566
rect 112 742 146 758
rect 112 550 146 566
rect -100 473 -84 507
rect 84 473 100 507
rect -100 365 -84 399
rect 84 365 100 399
rect -146 306 -112 322
rect -146 114 -112 130
rect 112 306 146 322
rect 112 114 146 130
rect -100 37 -84 71
rect 84 37 100 71
rect -100 -71 -84 -37
rect 84 -71 100 -37
rect -146 -130 -112 -114
rect -146 -322 -112 -306
rect 112 -130 146 -114
rect 112 -322 146 -306
rect -100 -399 -84 -365
rect 84 -399 100 -365
rect -100 -507 -84 -473
rect 84 -507 100 -473
rect -146 -566 -112 -550
rect -146 -758 -112 -742
rect 112 -566 146 -550
rect 112 -758 146 -742
rect -100 -835 -84 -801
rect 84 -835 100 -801
rect -100 -943 -84 -909
rect 84 -943 100 -909
rect -146 -1002 -112 -986
rect -146 -1194 -112 -1178
rect 112 -1002 146 -986
rect 112 -1194 146 -1178
rect -100 -1271 -84 -1237
rect 84 -1271 100 -1237
rect -100 -1379 -84 -1345
rect 84 -1379 100 -1345
rect -146 -1438 -112 -1422
rect -146 -1630 -112 -1614
rect 112 -1438 146 -1422
rect 112 -1630 146 -1614
rect -100 -1707 -84 -1673
rect 84 -1707 100 -1673
rect -100 -1815 -84 -1781
rect 84 -1815 100 -1781
rect -146 -1874 -112 -1858
rect -146 -2066 -112 -2050
rect 112 -1874 146 -1858
rect 112 -2066 146 -2050
rect -100 -2143 -84 -2109
rect 84 -2143 100 -2109
rect -100 -2251 -84 -2217
rect 84 -2251 100 -2217
rect -146 -2310 -112 -2294
rect -146 -2502 -112 -2486
rect 112 -2310 146 -2294
rect 112 -2502 146 -2486
rect -100 -2579 -84 -2545
rect 84 -2579 100 -2545
rect -100 -2687 -84 -2653
rect 84 -2687 100 -2653
rect -146 -2746 -112 -2730
rect -146 -2938 -112 -2922
rect 112 -2746 146 -2730
rect 112 -2938 146 -2922
rect -100 -3015 -84 -2981
rect 84 -3015 100 -2981
rect -100 -3123 -84 -3089
rect 84 -3123 100 -3089
rect -146 -3182 -112 -3166
rect -146 -3374 -112 -3358
rect 112 -3182 146 -3166
rect 112 -3374 146 -3358
rect -100 -3451 -84 -3417
rect 84 -3451 100 -3417
rect -100 -3559 -84 -3525
rect 84 -3559 100 -3525
rect -146 -3618 -112 -3602
rect -146 -3810 -112 -3794
rect 112 -3618 146 -3602
rect 112 -3810 146 -3794
rect -100 -3887 -84 -3853
rect 84 -3887 100 -3853
rect -100 -3995 -84 -3961
rect 84 -3995 100 -3961
rect -146 -4054 -112 -4038
rect -146 -4246 -112 -4230
rect 112 -4054 146 -4038
rect 112 -4246 146 -4230
rect -100 -4323 -84 -4289
rect 84 -4323 100 -4289
rect -100 -4431 -84 -4397
rect 84 -4431 100 -4397
rect -146 -4490 -112 -4474
rect -146 -4682 -112 -4666
rect 112 -4490 146 -4474
rect 112 -4682 146 -4666
rect -100 -4759 -84 -4725
rect 84 -4759 100 -4725
rect -100 -4867 -84 -4833
rect 84 -4867 100 -4833
rect -146 -4926 -112 -4910
rect -146 -5118 -112 -5102
rect 112 -4926 146 -4910
rect 112 -5118 146 -5102
rect -100 -5195 -84 -5161
rect 84 -5195 100 -5161
rect -100 -5303 -84 -5269
rect 84 -5303 100 -5269
rect -146 -5362 -112 -5346
rect -146 -5554 -112 -5538
rect 112 -5362 146 -5346
rect 112 -5554 146 -5538
rect -100 -5631 -84 -5597
rect 84 -5631 100 -5597
rect -100 -5739 -84 -5705
rect 84 -5739 100 -5705
rect -146 -5798 -112 -5782
rect -146 -5990 -112 -5974
rect 112 -5798 146 -5782
rect 112 -5990 146 -5974
rect -100 -6067 -84 -6033
rect 84 -6067 100 -6033
rect -260 -6135 -226 -6073
rect 226 -6135 260 -6073
rect -260 -6169 -164 -6135
rect 164 -6169 260 -6135
<< viali >>
rect -84 6033 84 6067
rect -146 5798 -112 5974
rect 112 5798 146 5974
rect -84 5705 84 5739
rect -84 5597 84 5631
rect -146 5362 -112 5538
rect 112 5362 146 5538
rect -84 5269 84 5303
rect -84 5161 84 5195
rect -146 4926 -112 5102
rect 112 4926 146 5102
rect -84 4833 84 4867
rect -84 4725 84 4759
rect -146 4490 -112 4666
rect 112 4490 146 4666
rect -84 4397 84 4431
rect -84 4289 84 4323
rect -146 4054 -112 4230
rect 112 4054 146 4230
rect -84 3961 84 3995
rect -84 3853 84 3887
rect -146 3618 -112 3794
rect 112 3618 146 3794
rect -84 3525 84 3559
rect -84 3417 84 3451
rect -146 3182 -112 3358
rect 112 3182 146 3358
rect -84 3089 84 3123
rect -84 2981 84 3015
rect -146 2746 -112 2922
rect 112 2746 146 2922
rect -84 2653 84 2687
rect -84 2545 84 2579
rect -146 2310 -112 2486
rect 112 2310 146 2486
rect -84 2217 84 2251
rect -84 2109 84 2143
rect -146 1874 -112 2050
rect 112 1874 146 2050
rect -84 1781 84 1815
rect -84 1673 84 1707
rect -146 1438 -112 1614
rect 112 1438 146 1614
rect -84 1345 84 1379
rect -84 1237 84 1271
rect -146 1002 -112 1178
rect 112 1002 146 1178
rect -84 909 84 943
rect -84 801 84 835
rect -146 566 -112 742
rect 112 566 146 742
rect -84 473 84 507
rect -84 365 84 399
rect -146 130 -112 306
rect 112 130 146 306
rect -84 37 84 71
rect -84 -71 84 -37
rect -146 -306 -112 -130
rect 112 -306 146 -130
rect -84 -399 84 -365
rect -84 -507 84 -473
rect -146 -742 -112 -566
rect 112 -742 146 -566
rect -84 -835 84 -801
rect -84 -943 84 -909
rect -146 -1178 -112 -1002
rect 112 -1178 146 -1002
rect -84 -1271 84 -1237
rect -84 -1379 84 -1345
rect -146 -1614 -112 -1438
rect 112 -1614 146 -1438
rect -84 -1707 84 -1673
rect -84 -1815 84 -1781
rect -146 -2050 -112 -1874
rect 112 -2050 146 -1874
rect -84 -2143 84 -2109
rect -84 -2251 84 -2217
rect -146 -2486 -112 -2310
rect 112 -2486 146 -2310
rect -84 -2579 84 -2545
rect -84 -2687 84 -2653
rect -146 -2922 -112 -2746
rect 112 -2922 146 -2746
rect -84 -3015 84 -2981
rect -84 -3123 84 -3089
rect -146 -3358 -112 -3182
rect 112 -3358 146 -3182
rect -84 -3451 84 -3417
rect -84 -3559 84 -3525
rect -146 -3794 -112 -3618
rect 112 -3794 146 -3618
rect -84 -3887 84 -3853
rect -84 -3995 84 -3961
rect -146 -4230 -112 -4054
rect 112 -4230 146 -4054
rect -84 -4323 84 -4289
rect -84 -4431 84 -4397
rect -146 -4666 -112 -4490
rect 112 -4666 146 -4490
rect -84 -4759 84 -4725
rect -84 -4867 84 -4833
rect -146 -5102 -112 -4926
rect 112 -5102 146 -4926
rect -84 -5195 84 -5161
rect -84 -5303 84 -5269
rect -146 -5538 -112 -5362
rect 112 -5538 146 -5362
rect -84 -5631 84 -5597
rect -84 -5739 84 -5705
rect -146 -5974 -112 -5798
rect 112 -5974 146 -5798
rect -84 -6067 84 -6033
<< metal1 >>
rect -96 6067 96 6073
rect -96 6033 -84 6067
rect 84 6033 96 6067
rect -96 6027 96 6033
rect -152 5974 -106 5986
rect -152 5798 -146 5974
rect -112 5798 -106 5974
rect -152 5786 -106 5798
rect 106 5974 152 5986
rect 106 5798 112 5974
rect 146 5798 152 5974
rect 106 5786 152 5798
rect -96 5739 96 5745
rect -96 5705 -84 5739
rect 84 5705 96 5739
rect -96 5699 96 5705
rect -96 5631 96 5637
rect -96 5597 -84 5631
rect 84 5597 96 5631
rect -96 5591 96 5597
rect -152 5538 -106 5550
rect -152 5362 -146 5538
rect -112 5362 -106 5538
rect -152 5350 -106 5362
rect 106 5538 152 5550
rect 106 5362 112 5538
rect 146 5362 152 5538
rect 106 5350 152 5362
rect -96 5303 96 5309
rect -96 5269 -84 5303
rect 84 5269 96 5303
rect -96 5263 96 5269
rect -96 5195 96 5201
rect -96 5161 -84 5195
rect 84 5161 96 5195
rect -96 5155 96 5161
rect -152 5102 -106 5114
rect -152 4926 -146 5102
rect -112 4926 -106 5102
rect -152 4914 -106 4926
rect 106 5102 152 5114
rect 106 4926 112 5102
rect 146 4926 152 5102
rect 106 4914 152 4926
rect -96 4867 96 4873
rect -96 4833 -84 4867
rect 84 4833 96 4867
rect -96 4827 96 4833
rect -96 4759 96 4765
rect -96 4725 -84 4759
rect 84 4725 96 4759
rect -96 4719 96 4725
rect -152 4666 -106 4678
rect -152 4490 -146 4666
rect -112 4490 -106 4666
rect -152 4478 -106 4490
rect 106 4666 152 4678
rect 106 4490 112 4666
rect 146 4490 152 4666
rect 106 4478 152 4490
rect -96 4431 96 4437
rect -96 4397 -84 4431
rect 84 4397 96 4431
rect -96 4391 96 4397
rect -96 4323 96 4329
rect -96 4289 -84 4323
rect 84 4289 96 4323
rect -96 4283 96 4289
rect -152 4230 -106 4242
rect -152 4054 -146 4230
rect -112 4054 -106 4230
rect -152 4042 -106 4054
rect 106 4230 152 4242
rect 106 4054 112 4230
rect 146 4054 152 4230
rect 106 4042 152 4054
rect -96 3995 96 4001
rect -96 3961 -84 3995
rect 84 3961 96 3995
rect -96 3955 96 3961
rect -96 3887 96 3893
rect -96 3853 -84 3887
rect 84 3853 96 3887
rect -96 3847 96 3853
rect -152 3794 -106 3806
rect -152 3618 -146 3794
rect -112 3618 -106 3794
rect -152 3606 -106 3618
rect 106 3794 152 3806
rect 106 3618 112 3794
rect 146 3618 152 3794
rect 106 3606 152 3618
rect -96 3559 96 3565
rect -96 3525 -84 3559
rect 84 3525 96 3559
rect -96 3519 96 3525
rect -96 3451 96 3457
rect -96 3417 -84 3451
rect 84 3417 96 3451
rect -96 3411 96 3417
rect -152 3358 -106 3370
rect -152 3182 -146 3358
rect -112 3182 -106 3358
rect -152 3170 -106 3182
rect 106 3358 152 3370
rect 106 3182 112 3358
rect 146 3182 152 3358
rect 106 3170 152 3182
rect -96 3123 96 3129
rect -96 3089 -84 3123
rect 84 3089 96 3123
rect -96 3083 96 3089
rect -96 3015 96 3021
rect -96 2981 -84 3015
rect 84 2981 96 3015
rect -96 2975 96 2981
rect -152 2922 -106 2934
rect -152 2746 -146 2922
rect -112 2746 -106 2922
rect -152 2734 -106 2746
rect 106 2922 152 2934
rect 106 2746 112 2922
rect 146 2746 152 2922
rect 106 2734 152 2746
rect -96 2687 96 2693
rect -96 2653 -84 2687
rect 84 2653 96 2687
rect -96 2647 96 2653
rect -96 2579 96 2585
rect -96 2545 -84 2579
rect 84 2545 96 2579
rect -96 2539 96 2545
rect -152 2486 -106 2498
rect -152 2310 -146 2486
rect -112 2310 -106 2486
rect -152 2298 -106 2310
rect 106 2486 152 2498
rect 106 2310 112 2486
rect 146 2310 152 2486
rect 106 2298 152 2310
rect -96 2251 96 2257
rect -96 2217 -84 2251
rect 84 2217 96 2251
rect -96 2211 96 2217
rect -96 2143 96 2149
rect -96 2109 -84 2143
rect 84 2109 96 2143
rect -96 2103 96 2109
rect -152 2050 -106 2062
rect -152 1874 -146 2050
rect -112 1874 -106 2050
rect -152 1862 -106 1874
rect 106 2050 152 2062
rect 106 1874 112 2050
rect 146 1874 152 2050
rect 106 1862 152 1874
rect -96 1815 96 1821
rect -96 1781 -84 1815
rect 84 1781 96 1815
rect -96 1775 96 1781
rect -96 1707 96 1713
rect -96 1673 -84 1707
rect 84 1673 96 1707
rect -96 1667 96 1673
rect -152 1614 -106 1626
rect -152 1438 -146 1614
rect -112 1438 -106 1614
rect -152 1426 -106 1438
rect 106 1614 152 1626
rect 106 1438 112 1614
rect 146 1438 152 1614
rect 106 1426 152 1438
rect -96 1379 96 1385
rect -96 1345 -84 1379
rect 84 1345 96 1379
rect -96 1339 96 1345
rect -96 1271 96 1277
rect -96 1237 -84 1271
rect 84 1237 96 1271
rect -96 1231 96 1237
rect -152 1178 -106 1190
rect -152 1002 -146 1178
rect -112 1002 -106 1178
rect -152 990 -106 1002
rect 106 1178 152 1190
rect 106 1002 112 1178
rect 146 1002 152 1178
rect 106 990 152 1002
rect -96 943 96 949
rect -96 909 -84 943
rect 84 909 96 943
rect -96 903 96 909
rect -96 835 96 841
rect -96 801 -84 835
rect 84 801 96 835
rect -96 795 96 801
rect -152 742 -106 754
rect -152 566 -146 742
rect -112 566 -106 742
rect -152 554 -106 566
rect 106 742 152 754
rect 106 566 112 742
rect 146 566 152 742
rect 106 554 152 566
rect -96 507 96 513
rect -96 473 -84 507
rect 84 473 96 507
rect -96 467 96 473
rect -96 399 96 405
rect -96 365 -84 399
rect 84 365 96 399
rect -96 359 96 365
rect -152 306 -106 318
rect -152 130 -146 306
rect -112 130 -106 306
rect -152 118 -106 130
rect 106 306 152 318
rect 106 130 112 306
rect 146 130 152 306
rect 106 118 152 130
rect -96 71 96 77
rect -96 37 -84 71
rect 84 37 96 71
rect -96 31 96 37
rect -96 -37 96 -31
rect -96 -71 -84 -37
rect 84 -71 96 -37
rect -96 -77 96 -71
rect -152 -130 -106 -118
rect -152 -306 -146 -130
rect -112 -306 -106 -130
rect -152 -318 -106 -306
rect 106 -130 152 -118
rect 106 -306 112 -130
rect 146 -306 152 -130
rect 106 -318 152 -306
rect -96 -365 96 -359
rect -96 -399 -84 -365
rect 84 -399 96 -365
rect -96 -405 96 -399
rect -96 -473 96 -467
rect -96 -507 -84 -473
rect 84 -507 96 -473
rect -96 -513 96 -507
rect -152 -566 -106 -554
rect -152 -742 -146 -566
rect -112 -742 -106 -566
rect -152 -754 -106 -742
rect 106 -566 152 -554
rect 106 -742 112 -566
rect 146 -742 152 -566
rect 106 -754 152 -742
rect -96 -801 96 -795
rect -96 -835 -84 -801
rect 84 -835 96 -801
rect -96 -841 96 -835
rect -96 -909 96 -903
rect -96 -943 -84 -909
rect 84 -943 96 -909
rect -96 -949 96 -943
rect -152 -1002 -106 -990
rect -152 -1178 -146 -1002
rect -112 -1178 -106 -1002
rect -152 -1190 -106 -1178
rect 106 -1002 152 -990
rect 106 -1178 112 -1002
rect 146 -1178 152 -1002
rect 106 -1190 152 -1178
rect -96 -1237 96 -1231
rect -96 -1271 -84 -1237
rect 84 -1271 96 -1237
rect -96 -1277 96 -1271
rect -96 -1345 96 -1339
rect -96 -1379 -84 -1345
rect 84 -1379 96 -1345
rect -96 -1385 96 -1379
rect -152 -1438 -106 -1426
rect -152 -1614 -146 -1438
rect -112 -1614 -106 -1438
rect -152 -1626 -106 -1614
rect 106 -1438 152 -1426
rect 106 -1614 112 -1438
rect 146 -1614 152 -1438
rect 106 -1626 152 -1614
rect -96 -1673 96 -1667
rect -96 -1707 -84 -1673
rect 84 -1707 96 -1673
rect -96 -1713 96 -1707
rect -96 -1781 96 -1775
rect -96 -1815 -84 -1781
rect 84 -1815 96 -1781
rect -96 -1821 96 -1815
rect -152 -1874 -106 -1862
rect -152 -2050 -146 -1874
rect -112 -2050 -106 -1874
rect -152 -2062 -106 -2050
rect 106 -1874 152 -1862
rect 106 -2050 112 -1874
rect 146 -2050 152 -1874
rect 106 -2062 152 -2050
rect -96 -2109 96 -2103
rect -96 -2143 -84 -2109
rect 84 -2143 96 -2109
rect -96 -2149 96 -2143
rect -96 -2217 96 -2211
rect -96 -2251 -84 -2217
rect 84 -2251 96 -2217
rect -96 -2257 96 -2251
rect -152 -2310 -106 -2298
rect -152 -2486 -146 -2310
rect -112 -2486 -106 -2310
rect -152 -2498 -106 -2486
rect 106 -2310 152 -2298
rect 106 -2486 112 -2310
rect 146 -2486 152 -2310
rect 106 -2498 152 -2486
rect -96 -2545 96 -2539
rect -96 -2579 -84 -2545
rect 84 -2579 96 -2545
rect -96 -2585 96 -2579
rect -96 -2653 96 -2647
rect -96 -2687 -84 -2653
rect 84 -2687 96 -2653
rect -96 -2693 96 -2687
rect -152 -2746 -106 -2734
rect -152 -2922 -146 -2746
rect -112 -2922 -106 -2746
rect -152 -2934 -106 -2922
rect 106 -2746 152 -2734
rect 106 -2922 112 -2746
rect 146 -2922 152 -2746
rect 106 -2934 152 -2922
rect -96 -2981 96 -2975
rect -96 -3015 -84 -2981
rect 84 -3015 96 -2981
rect -96 -3021 96 -3015
rect -96 -3089 96 -3083
rect -96 -3123 -84 -3089
rect 84 -3123 96 -3089
rect -96 -3129 96 -3123
rect -152 -3182 -106 -3170
rect -152 -3358 -146 -3182
rect -112 -3358 -106 -3182
rect -152 -3370 -106 -3358
rect 106 -3182 152 -3170
rect 106 -3358 112 -3182
rect 146 -3358 152 -3182
rect 106 -3370 152 -3358
rect -96 -3417 96 -3411
rect -96 -3451 -84 -3417
rect 84 -3451 96 -3417
rect -96 -3457 96 -3451
rect -96 -3525 96 -3519
rect -96 -3559 -84 -3525
rect 84 -3559 96 -3525
rect -96 -3565 96 -3559
rect -152 -3618 -106 -3606
rect -152 -3794 -146 -3618
rect -112 -3794 -106 -3618
rect -152 -3806 -106 -3794
rect 106 -3618 152 -3606
rect 106 -3794 112 -3618
rect 146 -3794 152 -3618
rect 106 -3806 152 -3794
rect -96 -3853 96 -3847
rect -96 -3887 -84 -3853
rect 84 -3887 96 -3853
rect -96 -3893 96 -3887
rect -96 -3961 96 -3955
rect -96 -3995 -84 -3961
rect 84 -3995 96 -3961
rect -96 -4001 96 -3995
rect -152 -4054 -106 -4042
rect -152 -4230 -146 -4054
rect -112 -4230 -106 -4054
rect -152 -4242 -106 -4230
rect 106 -4054 152 -4042
rect 106 -4230 112 -4054
rect 146 -4230 152 -4054
rect 106 -4242 152 -4230
rect -96 -4289 96 -4283
rect -96 -4323 -84 -4289
rect 84 -4323 96 -4289
rect -96 -4329 96 -4323
rect -96 -4397 96 -4391
rect -96 -4431 -84 -4397
rect 84 -4431 96 -4397
rect -96 -4437 96 -4431
rect -152 -4490 -106 -4478
rect -152 -4666 -146 -4490
rect -112 -4666 -106 -4490
rect -152 -4678 -106 -4666
rect 106 -4490 152 -4478
rect 106 -4666 112 -4490
rect 146 -4666 152 -4490
rect 106 -4678 152 -4666
rect -96 -4725 96 -4719
rect -96 -4759 -84 -4725
rect 84 -4759 96 -4725
rect -96 -4765 96 -4759
rect -96 -4833 96 -4827
rect -96 -4867 -84 -4833
rect 84 -4867 96 -4833
rect -96 -4873 96 -4867
rect -152 -4926 -106 -4914
rect -152 -5102 -146 -4926
rect -112 -5102 -106 -4926
rect -152 -5114 -106 -5102
rect 106 -4926 152 -4914
rect 106 -5102 112 -4926
rect 146 -5102 152 -4926
rect 106 -5114 152 -5102
rect -96 -5161 96 -5155
rect -96 -5195 -84 -5161
rect 84 -5195 96 -5161
rect -96 -5201 96 -5195
rect -96 -5269 96 -5263
rect -96 -5303 -84 -5269
rect 84 -5303 96 -5269
rect -96 -5309 96 -5303
rect -152 -5362 -106 -5350
rect -152 -5538 -146 -5362
rect -112 -5538 -106 -5362
rect -152 -5550 -106 -5538
rect 106 -5362 152 -5350
rect 106 -5538 112 -5362
rect 146 -5538 152 -5362
rect 106 -5550 152 -5538
rect -96 -5597 96 -5591
rect -96 -5631 -84 -5597
rect 84 -5631 96 -5597
rect -96 -5637 96 -5631
rect -96 -5705 96 -5699
rect -96 -5739 -84 -5705
rect 84 -5739 96 -5705
rect -96 -5745 96 -5739
rect -152 -5798 -106 -5786
rect -152 -5974 -146 -5798
rect -112 -5974 -106 -5798
rect -152 -5986 -106 -5974
rect 106 -5798 152 -5786
rect 106 -5974 112 -5798
rect 146 -5974 152 -5798
rect 106 -5986 152 -5974
rect -96 -6033 96 -6027
rect -96 -6067 -84 -6033
rect 84 -6067 96 -6033
rect -96 -6073 96 -6067
<< properties >>
string FIXED_BBOX -243 -6152 243 6152
string gencell sky130_fd_pr__pfet_01v8_lvt
string library sky130
string parameters w 1.0 l 1.0 m 28 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.35 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
