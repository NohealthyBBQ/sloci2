magic
tech sky130A
magscale 1 2
timestamp 1672437577
<< error_p >>
rect -2813 172 -2755 178
rect -2621 172 -2563 178
rect -2429 172 -2371 178
rect -2237 172 -2179 178
rect -2045 172 -1987 178
rect -1853 172 -1795 178
rect -1661 172 -1603 178
rect -1469 172 -1411 178
rect -1277 172 -1219 178
rect -1085 172 -1027 178
rect -893 172 -835 178
rect -701 172 -643 178
rect -509 172 -451 178
rect -317 172 -259 178
rect -125 172 -67 178
rect 67 172 125 178
rect 259 172 317 178
rect 451 172 509 178
rect 643 172 701 178
rect 835 172 893 178
rect 1027 172 1085 178
rect 1219 172 1277 178
rect 1411 172 1469 178
rect 1603 172 1661 178
rect 1795 172 1853 178
rect 1987 172 2045 178
rect 2179 172 2237 178
rect 2371 172 2429 178
rect 2563 172 2621 178
rect 2755 172 2813 178
rect -2813 138 -2801 172
rect -2621 138 -2609 172
rect -2429 138 -2417 172
rect -2237 138 -2225 172
rect -2045 138 -2033 172
rect -1853 138 -1841 172
rect -1661 138 -1649 172
rect -1469 138 -1457 172
rect -1277 138 -1265 172
rect -1085 138 -1073 172
rect -893 138 -881 172
rect -701 138 -689 172
rect -509 138 -497 172
rect -317 138 -305 172
rect -125 138 -113 172
rect 67 138 79 172
rect 259 138 271 172
rect 451 138 463 172
rect 643 138 655 172
rect 835 138 847 172
rect 1027 138 1039 172
rect 1219 138 1231 172
rect 1411 138 1423 172
rect 1603 138 1615 172
rect 1795 138 1807 172
rect 1987 138 1999 172
rect 2179 138 2191 172
rect 2371 138 2383 172
rect 2563 138 2575 172
rect 2755 138 2767 172
rect -2813 132 -2755 138
rect -2621 132 -2563 138
rect -2429 132 -2371 138
rect -2237 132 -2179 138
rect -2045 132 -1987 138
rect -1853 132 -1795 138
rect -1661 132 -1603 138
rect -1469 132 -1411 138
rect -1277 132 -1219 138
rect -1085 132 -1027 138
rect -893 132 -835 138
rect -701 132 -643 138
rect -509 132 -451 138
rect -317 132 -259 138
rect -125 132 -67 138
rect 67 132 125 138
rect 259 132 317 138
rect 451 132 509 138
rect 643 132 701 138
rect 835 132 893 138
rect 1027 132 1085 138
rect 1219 132 1277 138
rect 1411 132 1469 138
rect 1603 132 1661 138
rect 1795 132 1853 138
rect 1987 132 2045 138
rect 2179 132 2237 138
rect 2371 132 2429 138
rect 2563 132 2621 138
rect 2755 132 2813 138
rect -2909 -138 -2851 -132
rect -2717 -138 -2659 -132
rect -2525 -138 -2467 -132
rect -2333 -138 -2275 -132
rect -2141 -138 -2083 -132
rect -1949 -138 -1891 -132
rect -1757 -138 -1699 -132
rect -1565 -138 -1507 -132
rect -1373 -138 -1315 -132
rect -1181 -138 -1123 -132
rect -989 -138 -931 -132
rect -797 -138 -739 -132
rect -605 -138 -547 -132
rect -413 -138 -355 -132
rect -221 -138 -163 -132
rect -29 -138 29 -132
rect 163 -138 221 -132
rect 355 -138 413 -132
rect 547 -138 605 -132
rect 739 -138 797 -132
rect 931 -138 989 -132
rect 1123 -138 1181 -132
rect 1315 -138 1373 -132
rect 1507 -138 1565 -132
rect 1699 -138 1757 -132
rect 1891 -138 1949 -132
rect 2083 -138 2141 -132
rect 2275 -138 2333 -132
rect 2467 -138 2525 -132
rect 2659 -138 2717 -132
rect 2851 -138 2909 -132
rect -2909 -172 -2897 -138
rect -2717 -172 -2705 -138
rect -2525 -172 -2513 -138
rect -2333 -172 -2321 -138
rect -2141 -172 -2129 -138
rect -1949 -172 -1937 -138
rect -1757 -172 -1745 -138
rect -1565 -172 -1553 -138
rect -1373 -172 -1361 -138
rect -1181 -172 -1169 -138
rect -989 -172 -977 -138
rect -797 -172 -785 -138
rect -605 -172 -593 -138
rect -413 -172 -401 -138
rect -221 -172 -209 -138
rect -29 -172 -17 -138
rect 163 -172 175 -138
rect 355 -172 367 -138
rect 547 -172 559 -138
rect 739 -172 751 -138
rect 931 -172 943 -138
rect 1123 -172 1135 -138
rect 1315 -172 1327 -138
rect 1507 -172 1519 -138
rect 1699 -172 1711 -138
rect 1891 -172 1903 -138
rect 2083 -172 2095 -138
rect 2275 -172 2287 -138
rect 2467 -172 2479 -138
rect 2659 -172 2671 -138
rect 2851 -172 2863 -138
rect -2909 -178 -2851 -172
rect -2717 -178 -2659 -172
rect -2525 -178 -2467 -172
rect -2333 -178 -2275 -172
rect -2141 -178 -2083 -172
rect -1949 -178 -1891 -172
rect -1757 -178 -1699 -172
rect -1565 -178 -1507 -172
rect -1373 -178 -1315 -172
rect -1181 -178 -1123 -172
rect -989 -178 -931 -172
rect -797 -178 -739 -172
rect -605 -178 -547 -172
rect -413 -178 -355 -172
rect -221 -178 -163 -172
rect -29 -178 29 -172
rect 163 -178 221 -172
rect 355 -178 413 -172
rect 547 -178 605 -172
rect 739 -178 797 -172
rect 931 -178 989 -172
rect 1123 -178 1181 -172
rect 1315 -178 1373 -172
rect 1507 -178 1565 -172
rect 1699 -178 1757 -172
rect 1891 -178 1949 -172
rect 2083 -178 2141 -172
rect 2275 -178 2333 -172
rect 2467 -178 2525 -172
rect 2659 -178 2717 -172
rect 2851 -178 2909 -172
<< nmoslvt >>
rect -2895 -100 -2865 100
rect -2799 -100 -2769 100
rect -2703 -100 -2673 100
rect -2607 -100 -2577 100
rect -2511 -100 -2481 100
rect -2415 -100 -2385 100
rect -2319 -100 -2289 100
rect -2223 -100 -2193 100
rect -2127 -100 -2097 100
rect -2031 -100 -2001 100
rect -1935 -100 -1905 100
rect -1839 -100 -1809 100
rect -1743 -100 -1713 100
rect -1647 -100 -1617 100
rect -1551 -100 -1521 100
rect -1455 -100 -1425 100
rect -1359 -100 -1329 100
rect -1263 -100 -1233 100
rect -1167 -100 -1137 100
rect -1071 -100 -1041 100
rect -975 -100 -945 100
rect -879 -100 -849 100
rect -783 -100 -753 100
rect -687 -100 -657 100
rect -591 -100 -561 100
rect -495 -100 -465 100
rect -399 -100 -369 100
rect -303 -100 -273 100
rect -207 -100 -177 100
rect -111 -100 -81 100
rect -15 -100 15 100
rect 81 -100 111 100
rect 177 -100 207 100
rect 273 -100 303 100
rect 369 -100 399 100
rect 465 -100 495 100
rect 561 -100 591 100
rect 657 -100 687 100
rect 753 -100 783 100
rect 849 -100 879 100
rect 945 -100 975 100
rect 1041 -100 1071 100
rect 1137 -100 1167 100
rect 1233 -100 1263 100
rect 1329 -100 1359 100
rect 1425 -100 1455 100
rect 1521 -100 1551 100
rect 1617 -100 1647 100
rect 1713 -100 1743 100
rect 1809 -100 1839 100
rect 1905 -100 1935 100
rect 2001 -100 2031 100
rect 2097 -100 2127 100
rect 2193 -100 2223 100
rect 2289 -100 2319 100
rect 2385 -100 2415 100
rect 2481 -100 2511 100
rect 2577 -100 2607 100
rect 2673 -100 2703 100
rect 2769 -100 2799 100
rect 2865 -100 2895 100
<< ndiff >>
rect -2957 88 -2895 100
rect -2957 -88 -2945 88
rect -2911 -88 -2895 88
rect -2957 -100 -2895 -88
rect -2865 88 -2799 100
rect -2865 -88 -2849 88
rect -2815 -88 -2799 88
rect -2865 -100 -2799 -88
rect -2769 88 -2703 100
rect -2769 -88 -2753 88
rect -2719 -88 -2703 88
rect -2769 -100 -2703 -88
rect -2673 88 -2607 100
rect -2673 -88 -2657 88
rect -2623 -88 -2607 88
rect -2673 -100 -2607 -88
rect -2577 88 -2511 100
rect -2577 -88 -2561 88
rect -2527 -88 -2511 88
rect -2577 -100 -2511 -88
rect -2481 88 -2415 100
rect -2481 -88 -2465 88
rect -2431 -88 -2415 88
rect -2481 -100 -2415 -88
rect -2385 88 -2319 100
rect -2385 -88 -2369 88
rect -2335 -88 -2319 88
rect -2385 -100 -2319 -88
rect -2289 88 -2223 100
rect -2289 -88 -2273 88
rect -2239 -88 -2223 88
rect -2289 -100 -2223 -88
rect -2193 88 -2127 100
rect -2193 -88 -2177 88
rect -2143 -88 -2127 88
rect -2193 -100 -2127 -88
rect -2097 88 -2031 100
rect -2097 -88 -2081 88
rect -2047 -88 -2031 88
rect -2097 -100 -2031 -88
rect -2001 88 -1935 100
rect -2001 -88 -1985 88
rect -1951 -88 -1935 88
rect -2001 -100 -1935 -88
rect -1905 88 -1839 100
rect -1905 -88 -1889 88
rect -1855 -88 -1839 88
rect -1905 -100 -1839 -88
rect -1809 88 -1743 100
rect -1809 -88 -1793 88
rect -1759 -88 -1743 88
rect -1809 -100 -1743 -88
rect -1713 88 -1647 100
rect -1713 -88 -1697 88
rect -1663 -88 -1647 88
rect -1713 -100 -1647 -88
rect -1617 88 -1551 100
rect -1617 -88 -1601 88
rect -1567 -88 -1551 88
rect -1617 -100 -1551 -88
rect -1521 88 -1455 100
rect -1521 -88 -1505 88
rect -1471 -88 -1455 88
rect -1521 -100 -1455 -88
rect -1425 88 -1359 100
rect -1425 -88 -1409 88
rect -1375 -88 -1359 88
rect -1425 -100 -1359 -88
rect -1329 88 -1263 100
rect -1329 -88 -1313 88
rect -1279 -88 -1263 88
rect -1329 -100 -1263 -88
rect -1233 88 -1167 100
rect -1233 -88 -1217 88
rect -1183 -88 -1167 88
rect -1233 -100 -1167 -88
rect -1137 88 -1071 100
rect -1137 -88 -1121 88
rect -1087 -88 -1071 88
rect -1137 -100 -1071 -88
rect -1041 88 -975 100
rect -1041 -88 -1025 88
rect -991 -88 -975 88
rect -1041 -100 -975 -88
rect -945 88 -879 100
rect -945 -88 -929 88
rect -895 -88 -879 88
rect -945 -100 -879 -88
rect -849 88 -783 100
rect -849 -88 -833 88
rect -799 -88 -783 88
rect -849 -100 -783 -88
rect -753 88 -687 100
rect -753 -88 -737 88
rect -703 -88 -687 88
rect -753 -100 -687 -88
rect -657 88 -591 100
rect -657 -88 -641 88
rect -607 -88 -591 88
rect -657 -100 -591 -88
rect -561 88 -495 100
rect -561 -88 -545 88
rect -511 -88 -495 88
rect -561 -100 -495 -88
rect -465 88 -399 100
rect -465 -88 -449 88
rect -415 -88 -399 88
rect -465 -100 -399 -88
rect -369 88 -303 100
rect -369 -88 -353 88
rect -319 -88 -303 88
rect -369 -100 -303 -88
rect -273 88 -207 100
rect -273 -88 -257 88
rect -223 -88 -207 88
rect -273 -100 -207 -88
rect -177 88 -111 100
rect -177 -88 -161 88
rect -127 -88 -111 88
rect -177 -100 -111 -88
rect -81 88 -15 100
rect -81 -88 -65 88
rect -31 -88 -15 88
rect -81 -100 -15 -88
rect 15 88 81 100
rect 15 -88 31 88
rect 65 -88 81 88
rect 15 -100 81 -88
rect 111 88 177 100
rect 111 -88 127 88
rect 161 -88 177 88
rect 111 -100 177 -88
rect 207 88 273 100
rect 207 -88 223 88
rect 257 -88 273 88
rect 207 -100 273 -88
rect 303 88 369 100
rect 303 -88 319 88
rect 353 -88 369 88
rect 303 -100 369 -88
rect 399 88 465 100
rect 399 -88 415 88
rect 449 -88 465 88
rect 399 -100 465 -88
rect 495 88 561 100
rect 495 -88 511 88
rect 545 -88 561 88
rect 495 -100 561 -88
rect 591 88 657 100
rect 591 -88 607 88
rect 641 -88 657 88
rect 591 -100 657 -88
rect 687 88 753 100
rect 687 -88 703 88
rect 737 -88 753 88
rect 687 -100 753 -88
rect 783 88 849 100
rect 783 -88 799 88
rect 833 -88 849 88
rect 783 -100 849 -88
rect 879 88 945 100
rect 879 -88 895 88
rect 929 -88 945 88
rect 879 -100 945 -88
rect 975 88 1041 100
rect 975 -88 991 88
rect 1025 -88 1041 88
rect 975 -100 1041 -88
rect 1071 88 1137 100
rect 1071 -88 1087 88
rect 1121 -88 1137 88
rect 1071 -100 1137 -88
rect 1167 88 1233 100
rect 1167 -88 1183 88
rect 1217 -88 1233 88
rect 1167 -100 1233 -88
rect 1263 88 1329 100
rect 1263 -88 1279 88
rect 1313 -88 1329 88
rect 1263 -100 1329 -88
rect 1359 88 1425 100
rect 1359 -88 1375 88
rect 1409 -88 1425 88
rect 1359 -100 1425 -88
rect 1455 88 1521 100
rect 1455 -88 1471 88
rect 1505 -88 1521 88
rect 1455 -100 1521 -88
rect 1551 88 1617 100
rect 1551 -88 1567 88
rect 1601 -88 1617 88
rect 1551 -100 1617 -88
rect 1647 88 1713 100
rect 1647 -88 1663 88
rect 1697 -88 1713 88
rect 1647 -100 1713 -88
rect 1743 88 1809 100
rect 1743 -88 1759 88
rect 1793 -88 1809 88
rect 1743 -100 1809 -88
rect 1839 88 1905 100
rect 1839 -88 1855 88
rect 1889 -88 1905 88
rect 1839 -100 1905 -88
rect 1935 88 2001 100
rect 1935 -88 1951 88
rect 1985 -88 2001 88
rect 1935 -100 2001 -88
rect 2031 88 2097 100
rect 2031 -88 2047 88
rect 2081 -88 2097 88
rect 2031 -100 2097 -88
rect 2127 88 2193 100
rect 2127 -88 2143 88
rect 2177 -88 2193 88
rect 2127 -100 2193 -88
rect 2223 88 2289 100
rect 2223 -88 2239 88
rect 2273 -88 2289 88
rect 2223 -100 2289 -88
rect 2319 88 2385 100
rect 2319 -88 2335 88
rect 2369 -88 2385 88
rect 2319 -100 2385 -88
rect 2415 88 2481 100
rect 2415 -88 2431 88
rect 2465 -88 2481 88
rect 2415 -100 2481 -88
rect 2511 88 2577 100
rect 2511 -88 2527 88
rect 2561 -88 2577 88
rect 2511 -100 2577 -88
rect 2607 88 2673 100
rect 2607 -88 2623 88
rect 2657 -88 2673 88
rect 2607 -100 2673 -88
rect 2703 88 2769 100
rect 2703 -88 2719 88
rect 2753 -88 2769 88
rect 2703 -100 2769 -88
rect 2799 88 2865 100
rect 2799 -88 2815 88
rect 2849 -88 2865 88
rect 2799 -100 2865 -88
rect 2895 88 2957 100
rect 2895 -88 2911 88
rect 2945 -88 2957 88
rect 2895 -100 2957 -88
<< ndiffc >>
rect -2945 -88 -2911 88
rect -2849 -88 -2815 88
rect -2753 -88 -2719 88
rect -2657 -88 -2623 88
rect -2561 -88 -2527 88
rect -2465 -88 -2431 88
rect -2369 -88 -2335 88
rect -2273 -88 -2239 88
rect -2177 -88 -2143 88
rect -2081 -88 -2047 88
rect -1985 -88 -1951 88
rect -1889 -88 -1855 88
rect -1793 -88 -1759 88
rect -1697 -88 -1663 88
rect -1601 -88 -1567 88
rect -1505 -88 -1471 88
rect -1409 -88 -1375 88
rect -1313 -88 -1279 88
rect -1217 -88 -1183 88
rect -1121 -88 -1087 88
rect -1025 -88 -991 88
rect -929 -88 -895 88
rect -833 -88 -799 88
rect -737 -88 -703 88
rect -641 -88 -607 88
rect -545 -88 -511 88
rect -449 -88 -415 88
rect -353 -88 -319 88
rect -257 -88 -223 88
rect -161 -88 -127 88
rect -65 -88 -31 88
rect 31 -88 65 88
rect 127 -88 161 88
rect 223 -88 257 88
rect 319 -88 353 88
rect 415 -88 449 88
rect 511 -88 545 88
rect 607 -88 641 88
rect 703 -88 737 88
rect 799 -88 833 88
rect 895 -88 929 88
rect 991 -88 1025 88
rect 1087 -88 1121 88
rect 1183 -88 1217 88
rect 1279 -88 1313 88
rect 1375 -88 1409 88
rect 1471 -88 1505 88
rect 1567 -88 1601 88
rect 1663 -88 1697 88
rect 1759 -88 1793 88
rect 1855 -88 1889 88
rect 1951 -88 1985 88
rect 2047 -88 2081 88
rect 2143 -88 2177 88
rect 2239 -88 2273 88
rect 2335 -88 2369 88
rect 2431 -88 2465 88
rect 2527 -88 2561 88
rect 2623 -88 2657 88
rect 2719 -88 2753 88
rect 2815 -88 2849 88
rect 2911 -88 2945 88
<< poly >>
rect -2817 172 -2751 188
rect -2817 138 -2801 172
rect -2767 138 -2751 172
rect -2895 100 -2865 126
rect -2817 122 -2751 138
rect -2625 172 -2559 188
rect -2625 138 -2609 172
rect -2575 138 -2559 172
rect -2799 100 -2769 122
rect -2703 100 -2673 126
rect -2625 122 -2559 138
rect -2433 172 -2367 188
rect -2433 138 -2417 172
rect -2383 138 -2367 172
rect -2607 100 -2577 122
rect -2511 100 -2481 126
rect -2433 122 -2367 138
rect -2241 172 -2175 188
rect -2241 138 -2225 172
rect -2191 138 -2175 172
rect -2415 100 -2385 122
rect -2319 100 -2289 126
rect -2241 122 -2175 138
rect -2049 172 -1983 188
rect -2049 138 -2033 172
rect -1999 138 -1983 172
rect -2223 100 -2193 122
rect -2127 100 -2097 126
rect -2049 122 -1983 138
rect -1857 172 -1791 188
rect -1857 138 -1841 172
rect -1807 138 -1791 172
rect -2031 100 -2001 122
rect -1935 100 -1905 126
rect -1857 122 -1791 138
rect -1665 172 -1599 188
rect -1665 138 -1649 172
rect -1615 138 -1599 172
rect -1839 100 -1809 122
rect -1743 100 -1713 126
rect -1665 122 -1599 138
rect -1473 172 -1407 188
rect -1473 138 -1457 172
rect -1423 138 -1407 172
rect -1647 100 -1617 122
rect -1551 100 -1521 126
rect -1473 122 -1407 138
rect -1281 172 -1215 188
rect -1281 138 -1265 172
rect -1231 138 -1215 172
rect -1455 100 -1425 122
rect -1359 100 -1329 126
rect -1281 122 -1215 138
rect -1089 172 -1023 188
rect -1089 138 -1073 172
rect -1039 138 -1023 172
rect -1263 100 -1233 122
rect -1167 100 -1137 126
rect -1089 122 -1023 138
rect -897 172 -831 188
rect -897 138 -881 172
rect -847 138 -831 172
rect -1071 100 -1041 122
rect -975 100 -945 126
rect -897 122 -831 138
rect -705 172 -639 188
rect -705 138 -689 172
rect -655 138 -639 172
rect -879 100 -849 122
rect -783 100 -753 126
rect -705 122 -639 138
rect -513 172 -447 188
rect -513 138 -497 172
rect -463 138 -447 172
rect -687 100 -657 122
rect -591 100 -561 126
rect -513 122 -447 138
rect -321 172 -255 188
rect -321 138 -305 172
rect -271 138 -255 172
rect -495 100 -465 122
rect -399 100 -369 126
rect -321 122 -255 138
rect -129 172 -63 188
rect -129 138 -113 172
rect -79 138 -63 172
rect -303 100 -273 122
rect -207 100 -177 126
rect -129 122 -63 138
rect 63 172 129 188
rect 63 138 79 172
rect 113 138 129 172
rect -111 100 -81 122
rect -15 100 15 126
rect 63 122 129 138
rect 255 172 321 188
rect 255 138 271 172
rect 305 138 321 172
rect 81 100 111 122
rect 177 100 207 126
rect 255 122 321 138
rect 447 172 513 188
rect 447 138 463 172
rect 497 138 513 172
rect 273 100 303 122
rect 369 100 399 126
rect 447 122 513 138
rect 639 172 705 188
rect 639 138 655 172
rect 689 138 705 172
rect 465 100 495 122
rect 561 100 591 126
rect 639 122 705 138
rect 831 172 897 188
rect 831 138 847 172
rect 881 138 897 172
rect 657 100 687 122
rect 753 100 783 126
rect 831 122 897 138
rect 1023 172 1089 188
rect 1023 138 1039 172
rect 1073 138 1089 172
rect 849 100 879 122
rect 945 100 975 126
rect 1023 122 1089 138
rect 1215 172 1281 188
rect 1215 138 1231 172
rect 1265 138 1281 172
rect 1041 100 1071 122
rect 1137 100 1167 126
rect 1215 122 1281 138
rect 1407 172 1473 188
rect 1407 138 1423 172
rect 1457 138 1473 172
rect 1233 100 1263 122
rect 1329 100 1359 126
rect 1407 122 1473 138
rect 1599 172 1665 188
rect 1599 138 1615 172
rect 1649 138 1665 172
rect 1425 100 1455 122
rect 1521 100 1551 126
rect 1599 122 1665 138
rect 1791 172 1857 188
rect 1791 138 1807 172
rect 1841 138 1857 172
rect 1617 100 1647 122
rect 1713 100 1743 126
rect 1791 122 1857 138
rect 1983 172 2049 188
rect 1983 138 1999 172
rect 2033 138 2049 172
rect 1809 100 1839 122
rect 1905 100 1935 126
rect 1983 122 2049 138
rect 2175 172 2241 188
rect 2175 138 2191 172
rect 2225 138 2241 172
rect 2001 100 2031 122
rect 2097 100 2127 126
rect 2175 122 2241 138
rect 2367 172 2433 188
rect 2367 138 2383 172
rect 2417 138 2433 172
rect 2193 100 2223 122
rect 2289 100 2319 126
rect 2367 122 2433 138
rect 2559 172 2625 188
rect 2559 138 2575 172
rect 2609 138 2625 172
rect 2385 100 2415 122
rect 2481 100 2511 126
rect 2559 122 2625 138
rect 2751 172 2817 188
rect 2751 138 2767 172
rect 2801 138 2817 172
rect 2577 100 2607 122
rect 2673 100 2703 126
rect 2751 122 2817 138
rect 2769 100 2799 122
rect 2865 100 2895 126
rect -2895 -122 -2865 -100
rect -2913 -138 -2847 -122
rect -2799 -126 -2769 -100
rect -2703 -122 -2673 -100
rect -2913 -172 -2897 -138
rect -2863 -172 -2847 -138
rect -2913 -188 -2847 -172
rect -2721 -138 -2655 -122
rect -2607 -126 -2577 -100
rect -2511 -122 -2481 -100
rect -2721 -172 -2705 -138
rect -2671 -172 -2655 -138
rect -2721 -188 -2655 -172
rect -2529 -138 -2463 -122
rect -2415 -126 -2385 -100
rect -2319 -122 -2289 -100
rect -2529 -172 -2513 -138
rect -2479 -172 -2463 -138
rect -2529 -188 -2463 -172
rect -2337 -138 -2271 -122
rect -2223 -126 -2193 -100
rect -2127 -122 -2097 -100
rect -2337 -172 -2321 -138
rect -2287 -172 -2271 -138
rect -2337 -188 -2271 -172
rect -2145 -138 -2079 -122
rect -2031 -126 -2001 -100
rect -1935 -122 -1905 -100
rect -2145 -172 -2129 -138
rect -2095 -172 -2079 -138
rect -2145 -188 -2079 -172
rect -1953 -138 -1887 -122
rect -1839 -126 -1809 -100
rect -1743 -122 -1713 -100
rect -1953 -172 -1937 -138
rect -1903 -172 -1887 -138
rect -1953 -188 -1887 -172
rect -1761 -138 -1695 -122
rect -1647 -126 -1617 -100
rect -1551 -122 -1521 -100
rect -1761 -172 -1745 -138
rect -1711 -172 -1695 -138
rect -1761 -188 -1695 -172
rect -1569 -138 -1503 -122
rect -1455 -126 -1425 -100
rect -1359 -122 -1329 -100
rect -1569 -172 -1553 -138
rect -1519 -172 -1503 -138
rect -1569 -188 -1503 -172
rect -1377 -138 -1311 -122
rect -1263 -126 -1233 -100
rect -1167 -122 -1137 -100
rect -1377 -172 -1361 -138
rect -1327 -172 -1311 -138
rect -1377 -188 -1311 -172
rect -1185 -138 -1119 -122
rect -1071 -126 -1041 -100
rect -975 -122 -945 -100
rect -1185 -172 -1169 -138
rect -1135 -172 -1119 -138
rect -1185 -188 -1119 -172
rect -993 -138 -927 -122
rect -879 -126 -849 -100
rect -783 -122 -753 -100
rect -993 -172 -977 -138
rect -943 -172 -927 -138
rect -993 -188 -927 -172
rect -801 -138 -735 -122
rect -687 -126 -657 -100
rect -591 -122 -561 -100
rect -801 -172 -785 -138
rect -751 -172 -735 -138
rect -801 -188 -735 -172
rect -609 -138 -543 -122
rect -495 -126 -465 -100
rect -399 -122 -369 -100
rect -609 -172 -593 -138
rect -559 -172 -543 -138
rect -609 -188 -543 -172
rect -417 -138 -351 -122
rect -303 -126 -273 -100
rect -207 -122 -177 -100
rect -417 -172 -401 -138
rect -367 -172 -351 -138
rect -417 -188 -351 -172
rect -225 -138 -159 -122
rect -111 -126 -81 -100
rect -15 -122 15 -100
rect -225 -172 -209 -138
rect -175 -172 -159 -138
rect -225 -188 -159 -172
rect -33 -138 33 -122
rect 81 -126 111 -100
rect 177 -122 207 -100
rect -33 -172 -17 -138
rect 17 -172 33 -138
rect -33 -188 33 -172
rect 159 -138 225 -122
rect 273 -126 303 -100
rect 369 -122 399 -100
rect 159 -172 175 -138
rect 209 -172 225 -138
rect 159 -188 225 -172
rect 351 -138 417 -122
rect 465 -126 495 -100
rect 561 -122 591 -100
rect 351 -172 367 -138
rect 401 -172 417 -138
rect 351 -188 417 -172
rect 543 -138 609 -122
rect 657 -126 687 -100
rect 753 -122 783 -100
rect 543 -172 559 -138
rect 593 -172 609 -138
rect 543 -188 609 -172
rect 735 -138 801 -122
rect 849 -126 879 -100
rect 945 -122 975 -100
rect 735 -172 751 -138
rect 785 -172 801 -138
rect 735 -188 801 -172
rect 927 -138 993 -122
rect 1041 -126 1071 -100
rect 1137 -122 1167 -100
rect 927 -172 943 -138
rect 977 -172 993 -138
rect 927 -188 993 -172
rect 1119 -138 1185 -122
rect 1233 -126 1263 -100
rect 1329 -122 1359 -100
rect 1119 -172 1135 -138
rect 1169 -172 1185 -138
rect 1119 -188 1185 -172
rect 1311 -138 1377 -122
rect 1425 -126 1455 -100
rect 1521 -122 1551 -100
rect 1311 -172 1327 -138
rect 1361 -172 1377 -138
rect 1311 -188 1377 -172
rect 1503 -138 1569 -122
rect 1617 -126 1647 -100
rect 1713 -122 1743 -100
rect 1503 -172 1519 -138
rect 1553 -172 1569 -138
rect 1503 -188 1569 -172
rect 1695 -138 1761 -122
rect 1809 -126 1839 -100
rect 1905 -122 1935 -100
rect 1695 -172 1711 -138
rect 1745 -172 1761 -138
rect 1695 -188 1761 -172
rect 1887 -138 1953 -122
rect 2001 -126 2031 -100
rect 2097 -122 2127 -100
rect 1887 -172 1903 -138
rect 1937 -172 1953 -138
rect 1887 -188 1953 -172
rect 2079 -138 2145 -122
rect 2193 -126 2223 -100
rect 2289 -122 2319 -100
rect 2079 -172 2095 -138
rect 2129 -172 2145 -138
rect 2079 -188 2145 -172
rect 2271 -138 2337 -122
rect 2385 -126 2415 -100
rect 2481 -122 2511 -100
rect 2271 -172 2287 -138
rect 2321 -172 2337 -138
rect 2271 -188 2337 -172
rect 2463 -138 2529 -122
rect 2577 -126 2607 -100
rect 2673 -122 2703 -100
rect 2463 -172 2479 -138
rect 2513 -172 2529 -138
rect 2463 -188 2529 -172
rect 2655 -138 2721 -122
rect 2769 -126 2799 -100
rect 2865 -122 2895 -100
rect 2655 -172 2671 -138
rect 2705 -172 2721 -138
rect 2655 -188 2721 -172
rect 2847 -138 2913 -122
rect 2847 -172 2863 -138
rect 2897 -172 2913 -138
rect 2847 -188 2913 -172
<< polycont >>
rect -2801 138 -2767 172
rect -2609 138 -2575 172
rect -2417 138 -2383 172
rect -2225 138 -2191 172
rect -2033 138 -1999 172
rect -1841 138 -1807 172
rect -1649 138 -1615 172
rect -1457 138 -1423 172
rect -1265 138 -1231 172
rect -1073 138 -1039 172
rect -881 138 -847 172
rect -689 138 -655 172
rect -497 138 -463 172
rect -305 138 -271 172
rect -113 138 -79 172
rect 79 138 113 172
rect 271 138 305 172
rect 463 138 497 172
rect 655 138 689 172
rect 847 138 881 172
rect 1039 138 1073 172
rect 1231 138 1265 172
rect 1423 138 1457 172
rect 1615 138 1649 172
rect 1807 138 1841 172
rect 1999 138 2033 172
rect 2191 138 2225 172
rect 2383 138 2417 172
rect 2575 138 2609 172
rect 2767 138 2801 172
rect -2897 -172 -2863 -138
rect -2705 -172 -2671 -138
rect -2513 -172 -2479 -138
rect -2321 -172 -2287 -138
rect -2129 -172 -2095 -138
rect -1937 -172 -1903 -138
rect -1745 -172 -1711 -138
rect -1553 -172 -1519 -138
rect -1361 -172 -1327 -138
rect -1169 -172 -1135 -138
rect -977 -172 -943 -138
rect -785 -172 -751 -138
rect -593 -172 -559 -138
rect -401 -172 -367 -138
rect -209 -172 -175 -138
rect -17 -172 17 -138
rect 175 -172 209 -138
rect 367 -172 401 -138
rect 559 -172 593 -138
rect 751 -172 785 -138
rect 943 -172 977 -138
rect 1135 -172 1169 -138
rect 1327 -172 1361 -138
rect 1519 -172 1553 -138
rect 1711 -172 1745 -138
rect 1903 -172 1937 -138
rect 2095 -172 2129 -138
rect 2287 -172 2321 -138
rect 2479 -172 2513 -138
rect 2671 -172 2705 -138
rect 2863 -172 2897 -138
<< locali >>
rect -2817 138 -2801 172
rect -2767 138 -2751 172
rect -2625 138 -2609 172
rect -2575 138 -2559 172
rect -2433 138 -2417 172
rect -2383 138 -2367 172
rect -2241 138 -2225 172
rect -2191 138 -2175 172
rect -2049 138 -2033 172
rect -1999 138 -1983 172
rect -1857 138 -1841 172
rect -1807 138 -1791 172
rect -1665 138 -1649 172
rect -1615 138 -1599 172
rect -1473 138 -1457 172
rect -1423 138 -1407 172
rect -1281 138 -1265 172
rect -1231 138 -1215 172
rect -1089 138 -1073 172
rect -1039 138 -1023 172
rect -897 138 -881 172
rect -847 138 -831 172
rect -705 138 -689 172
rect -655 138 -639 172
rect -513 138 -497 172
rect -463 138 -447 172
rect -321 138 -305 172
rect -271 138 -255 172
rect -129 138 -113 172
rect -79 138 -63 172
rect 63 138 79 172
rect 113 138 129 172
rect 255 138 271 172
rect 305 138 321 172
rect 447 138 463 172
rect 497 138 513 172
rect 639 138 655 172
rect 689 138 705 172
rect 831 138 847 172
rect 881 138 897 172
rect 1023 138 1039 172
rect 1073 138 1089 172
rect 1215 138 1231 172
rect 1265 138 1281 172
rect 1407 138 1423 172
rect 1457 138 1473 172
rect 1599 138 1615 172
rect 1649 138 1665 172
rect 1791 138 1807 172
rect 1841 138 1857 172
rect 1983 138 1999 172
rect 2033 138 2049 172
rect 2175 138 2191 172
rect 2225 138 2241 172
rect 2367 138 2383 172
rect 2417 138 2433 172
rect 2559 138 2575 172
rect 2609 138 2625 172
rect 2751 138 2767 172
rect 2801 138 2817 172
rect -2945 88 -2911 104
rect -2945 -104 -2911 -88
rect -2849 88 -2815 104
rect -2849 -104 -2815 -88
rect -2753 88 -2719 104
rect -2753 -104 -2719 -88
rect -2657 88 -2623 104
rect -2657 -104 -2623 -88
rect -2561 88 -2527 104
rect -2561 -104 -2527 -88
rect -2465 88 -2431 104
rect -2465 -104 -2431 -88
rect -2369 88 -2335 104
rect -2369 -104 -2335 -88
rect -2273 88 -2239 104
rect -2273 -104 -2239 -88
rect -2177 88 -2143 104
rect -2177 -104 -2143 -88
rect -2081 88 -2047 104
rect -2081 -104 -2047 -88
rect -1985 88 -1951 104
rect -1985 -104 -1951 -88
rect -1889 88 -1855 104
rect -1889 -104 -1855 -88
rect -1793 88 -1759 104
rect -1793 -104 -1759 -88
rect -1697 88 -1663 104
rect -1697 -104 -1663 -88
rect -1601 88 -1567 104
rect -1601 -104 -1567 -88
rect -1505 88 -1471 104
rect -1505 -104 -1471 -88
rect -1409 88 -1375 104
rect -1409 -104 -1375 -88
rect -1313 88 -1279 104
rect -1313 -104 -1279 -88
rect -1217 88 -1183 104
rect -1217 -104 -1183 -88
rect -1121 88 -1087 104
rect -1121 -104 -1087 -88
rect -1025 88 -991 104
rect -1025 -104 -991 -88
rect -929 88 -895 104
rect -929 -104 -895 -88
rect -833 88 -799 104
rect -833 -104 -799 -88
rect -737 88 -703 104
rect -737 -104 -703 -88
rect -641 88 -607 104
rect -641 -104 -607 -88
rect -545 88 -511 104
rect -545 -104 -511 -88
rect -449 88 -415 104
rect -449 -104 -415 -88
rect -353 88 -319 104
rect -353 -104 -319 -88
rect -257 88 -223 104
rect -257 -104 -223 -88
rect -161 88 -127 104
rect -161 -104 -127 -88
rect -65 88 -31 104
rect -65 -104 -31 -88
rect 31 88 65 104
rect 31 -104 65 -88
rect 127 88 161 104
rect 127 -104 161 -88
rect 223 88 257 104
rect 223 -104 257 -88
rect 319 88 353 104
rect 319 -104 353 -88
rect 415 88 449 104
rect 415 -104 449 -88
rect 511 88 545 104
rect 511 -104 545 -88
rect 607 88 641 104
rect 607 -104 641 -88
rect 703 88 737 104
rect 703 -104 737 -88
rect 799 88 833 104
rect 799 -104 833 -88
rect 895 88 929 104
rect 895 -104 929 -88
rect 991 88 1025 104
rect 991 -104 1025 -88
rect 1087 88 1121 104
rect 1087 -104 1121 -88
rect 1183 88 1217 104
rect 1183 -104 1217 -88
rect 1279 88 1313 104
rect 1279 -104 1313 -88
rect 1375 88 1409 104
rect 1375 -104 1409 -88
rect 1471 88 1505 104
rect 1471 -104 1505 -88
rect 1567 88 1601 104
rect 1567 -104 1601 -88
rect 1663 88 1697 104
rect 1663 -104 1697 -88
rect 1759 88 1793 104
rect 1759 -104 1793 -88
rect 1855 88 1889 104
rect 1855 -104 1889 -88
rect 1951 88 1985 104
rect 1951 -104 1985 -88
rect 2047 88 2081 104
rect 2047 -104 2081 -88
rect 2143 88 2177 104
rect 2143 -104 2177 -88
rect 2239 88 2273 104
rect 2239 -104 2273 -88
rect 2335 88 2369 104
rect 2335 -104 2369 -88
rect 2431 88 2465 104
rect 2431 -104 2465 -88
rect 2527 88 2561 104
rect 2527 -104 2561 -88
rect 2623 88 2657 104
rect 2623 -104 2657 -88
rect 2719 88 2753 104
rect 2719 -104 2753 -88
rect 2815 88 2849 104
rect 2815 -104 2849 -88
rect 2911 88 2945 104
rect 2911 -104 2945 -88
rect -2913 -172 -2897 -138
rect -2863 -172 -2847 -138
rect -2721 -172 -2705 -138
rect -2671 -172 -2655 -138
rect -2529 -172 -2513 -138
rect -2479 -172 -2463 -138
rect -2337 -172 -2321 -138
rect -2287 -172 -2271 -138
rect -2145 -172 -2129 -138
rect -2095 -172 -2079 -138
rect -1953 -172 -1937 -138
rect -1903 -172 -1887 -138
rect -1761 -172 -1745 -138
rect -1711 -172 -1695 -138
rect -1569 -172 -1553 -138
rect -1519 -172 -1503 -138
rect -1377 -172 -1361 -138
rect -1327 -172 -1311 -138
rect -1185 -172 -1169 -138
rect -1135 -172 -1119 -138
rect -993 -172 -977 -138
rect -943 -172 -927 -138
rect -801 -172 -785 -138
rect -751 -172 -735 -138
rect -609 -172 -593 -138
rect -559 -172 -543 -138
rect -417 -172 -401 -138
rect -367 -172 -351 -138
rect -225 -172 -209 -138
rect -175 -172 -159 -138
rect -33 -172 -17 -138
rect 17 -172 33 -138
rect 159 -172 175 -138
rect 209 -172 225 -138
rect 351 -172 367 -138
rect 401 -172 417 -138
rect 543 -172 559 -138
rect 593 -172 609 -138
rect 735 -172 751 -138
rect 785 -172 801 -138
rect 927 -172 943 -138
rect 977 -172 993 -138
rect 1119 -172 1135 -138
rect 1169 -172 1185 -138
rect 1311 -172 1327 -138
rect 1361 -172 1377 -138
rect 1503 -172 1519 -138
rect 1553 -172 1569 -138
rect 1695 -172 1711 -138
rect 1745 -172 1761 -138
rect 1887 -172 1903 -138
rect 1937 -172 1953 -138
rect 2079 -172 2095 -138
rect 2129 -172 2145 -138
rect 2271 -172 2287 -138
rect 2321 -172 2337 -138
rect 2463 -172 2479 -138
rect 2513 -172 2529 -138
rect 2655 -172 2671 -138
rect 2705 -172 2721 -138
rect 2847 -172 2863 -138
rect 2897 -172 2913 -138
<< viali >>
rect -2801 138 -2767 172
rect -2609 138 -2575 172
rect -2417 138 -2383 172
rect -2225 138 -2191 172
rect -2033 138 -1999 172
rect -1841 138 -1807 172
rect -1649 138 -1615 172
rect -1457 138 -1423 172
rect -1265 138 -1231 172
rect -1073 138 -1039 172
rect -881 138 -847 172
rect -689 138 -655 172
rect -497 138 -463 172
rect -305 138 -271 172
rect -113 138 -79 172
rect 79 138 113 172
rect 271 138 305 172
rect 463 138 497 172
rect 655 138 689 172
rect 847 138 881 172
rect 1039 138 1073 172
rect 1231 138 1265 172
rect 1423 138 1457 172
rect 1615 138 1649 172
rect 1807 138 1841 172
rect 1999 138 2033 172
rect 2191 138 2225 172
rect 2383 138 2417 172
rect 2575 138 2609 172
rect 2767 138 2801 172
rect -2945 -88 -2911 88
rect -2849 -88 -2815 88
rect -2753 -88 -2719 88
rect -2657 -88 -2623 88
rect -2561 -88 -2527 88
rect -2465 -88 -2431 88
rect -2369 -88 -2335 88
rect -2273 -88 -2239 88
rect -2177 -88 -2143 88
rect -2081 -88 -2047 88
rect -1985 -88 -1951 88
rect -1889 -88 -1855 88
rect -1793 -88 -1759 88
rect -1697 -88 -1663 88
rect -1601 -88 -1567 88
rect -1505 -88 -1471 88
rect -1409 -88 -1375 88
rect -1313 -88 -1279 88
rect -1217 -88 -1183 88
rect -1121 -88 -1087 88
rect -1025 -88 -991 88
rect -929 -88 -895 88
rect -833 -88 -799 88
rect -737 -88 -703 88
rect -641 -88 -607 88
rect -545 -88 -511 88
rect -449 -88 -415 88
rect -353 -88 -319 88
rect -257 -88 -223 88
rect -161 -88 -127 88
rect -65 -88 -31 88
rect 31 -88 65 88
rect 127 -88 161 88
rect 223 -88 257 88
rect 319 -88 353 88
rect 415 -88 449 88
rect 511 -88 545 88
rect 607 -88 641 88
rect 703 -88 737 88
rect 799 -88 833 88
rect 895 -88 929 88
rect 991 -88 1025 88
rect 1087 -88 1121 88
rect 1183 -88 1217 88
rect 1279 -88 1313 88
rect 1375 -88 1409 88
rect 1471 -88 1505 88
rect 1567 -88 1601 88
rect 1663 -88 1697 88
rect 1759 -88 1793 88
rect 1855 -88 1889 88
rect 1951 -88 1985 88
rect 2047 -88 2081 88
rect 2143 -88 2177 88
rect 2239 -88 2273 88
rect 2335 -88 2369 88
rect 2431 -88 2465 88
rect 2527 -88 2561 88
rect 2623 -88 2657 88
rect 2719 -88 2753 88
rect 2815 -88 2849 88
rect 2911 -88 2945 88
rect -2897 -172 -2863 -138
rect -2705 -172 -2671 -138
rect -2513 -172 -2479 -138
rect -2321 -172 -2287 -138
rect -2129 -172 -2095 -138
rect -1937 -172 -1903 -138
rect -1745 -172 -1711 -138
rect -1553 -172 -1519 -138
rect -1361 -172 -1327 -138
rect -1169 -172 -1135 -138
rect -977 -172 -943 -138
rect -785 -172 -751 -138
rect -593 -172 -559 -138
rect -401 -172 -367 -138
rect -209 -172 -175 -138
rect -17 -172 17 -138
rect 175 -172 209 -138
rect 367 -172 401 -138
rect 559 -172 593 -138
rect 751 -172 785 -138
rect 943 -172 977 -138
rect 1135 -172 1169 -138
rect 1327 -172 1361 -138
rect 1519 -172 1553 -138
rect 1711 -172 1745 -138
rect 1903 -172 1937 -138
rect 2095 -172 2129 -138
rect 2287 -172 2321 -138
rect 2479 -172 2513 -138
rect 2671 -172 2705 -138
rect 2863 -172 2897 -138
<< metal1 >>
rect -2813 172 -2755 178
rect -2813 138 -2801 172
rect -2767 138 -2755 172
rect -2813 132 -2755 138
rect -2621 172 -2563 178
rect -2621 138 -2609 172
rect -2575 138 -2563 172
rect -2621 132 -2563 138
rect -2429 172 -2371 178
rect -2429 138 -2417 172
rect -2383 138 -2371 172
rect -2429 132 -2371 138
rect -2237 172 -2179 178
rect -2237 138 -2225 172
rect -2191 138 -2179 172
rect -2237 132 -2179 138
rect -2045 172 -1987 178
rect -2045 138 -2033 172
rect -1999 138 -1987 172
rect -2045 132 -1987 138
rect -1853 172 -1795 178
rect -1853 138 -1841 172
rect -1807 138 -1795 172
rect -1853 132 -1795 138
rect -1661 172 -1603 178
rect -1661 138 -1649 172
rect -1615 138 -1603 172
rect -1661 132 -1603 138
rect -1469 172 -1411 178
rect -1469 138 -1457 172
rect -1423 138 -1411 172
rect -1469 132 -1411 138
rect -1277 172 -1219 178
rect -1277 138 -1265 172
rect -1231 138 -1219 172
rect -1277 132 -1219 138
rect -1085 172 -1027 178
rect -1085 138 -1073 172
rect -1039 138 -1027 172
rect -1085 132 -1027 138
rect -893 172 -835 178
rect -893 138 -881 172
rect -847 138 -835 172
rect -893 132 -835 138
rect -701 172 -643 178
rect -701 138 -689 172
rect -655 138 -643 172
rect -701 132 -643 138
rect -509 172 -451 178
rect -509 138 -497 172
rect -463 138 -451 172
rect -509 132 -451 138
rect -317 172 -259 178
rect -317 138 -305 172
rect -271 138 -259 172
rect -317 132 -259 138
rect -125 172 -67 178
rect -125 138 -113 172
rect -79 138 -67 172
rect -125 132 -67 138
rect 67 172 125 178
rect 67 138 79 172
rect 113 138 125 172
rect 67 132 125 138
rect 259 172 317 178
rect 259 138 271 172
rect 305 138 317 172
rect 259 132 317 138
rect 451 172 509 178
rect 451 138 463 172
rect 497 138 509 172
rect 451 132 509 138
rect 643 172 701 178
rect 643 138 655 172
rect 689 138 701 172
rect 643 132 701 138
rect 835 172 893 178
rect 835 138 847 172
rect 881 138 893 172
rect 835 132 893 138
rect 1027 172 1085 178
rect 1027 138 1039 172
rect 1073 138 1085 172
rect 1027 132 1085 138
rect 1219 172 1277 178
rect 1219 138 1231 172
rect 1265 138 1277 172
rect 1219 132 1277 138
rect 1411 172 1469 178
rect 1411 138 1423 172
rect 1457 138 1469 172
rect 1411 132 1469 138
rect 1603 172 1661 178
rect 1603 138 1615 172
rect 1649 138 1661 172
rect 1603 132 1661 138
rect 1795 172 1853 178
rect 1795 138 1807 172
rect 1841 138 1853 172
rect 1795 132 1853 138
rect 1987 172 2045 178
rect 1987 138 1999 172
rect 2033 138 2045 172
rect 1987 132 2045 138
rect 2179 172 2237 178
rect 2179 138 2191 172
rect 2225 138 2237 172
rect 2179 132 2237 138
rect 2371 172 2429 178
rect 2371 138 2383 172
rect 2417 138 2429 172
rect 2371 132 2429 138
rect 2563 172 2621 178
rect 2563 138 2575 172
rect 2609 138 2621 172
rect 2563 132 2621 138
rect 2755 172 2813 178
rect 2755 138 2767 172
rect 2801 138 2813 172
rect 2755 132 2813 138
rect -2951 88 -2905 100
rect -2951 -88 -2945 88
rect -2911 -88 -2905 88
rect -2951 -100 -2905 -88
rect -2855 88 -2809 100
rect -2855 -88 -2849 88
rect -2815 -88 -2809 88
rect -2855 -100 -2809 -88
rect -2759 88 -2713 100
rect -2759 -88 -2753 88
rect -2719 -88 -2713 88
rect -2759 -100 -2713 -88
rect -2663 88 -2617 100
rect -2663 -88 -2657 88
rect -2623 -88 -2617 88
rect -2663 -100 -2617 -88
rect -2567 88 -2521 100
rect -2567 -88 -2561 88
rect -2527 -88 -2521 88
rect -2567 -100 -2521 -88
rect -2471 88 -2425 100
rect -2471 -88 -2465 88
rect -2431 -88 -2425 88
rect -2471 -100 -2425 -88
rect -2375 88 -2329 100
rect -2375 -88 -2369 88
rect -2335 -88 -2329 88
rect -2375 -100 -2329 -88
rect -2279 88 -2233 100
rect -2279 -88 -2273 88
rect -2239 -88 -2233 88
rect -2279 -100 -2233 -88
rect -2183 88 -2137 100
rect -2183 -88 -2177 88
rect -2143 -88 -2137 88
rect -2183 -100 -2137 -88
rect -2087 88 -2041 100
rect -2087 -88 -2081 88
rect -2047 -88 -2041 88
rect -2087 -100 -2041 -88
rect -1991 88 -1945 100
rect -1991 -88 -1985 88
rect -1951 -88 -1945 88
rect -1991 -100 -1945 -88
rect -1895 88 -1849 100
rect -1895 -88 -1889 88
rect -1855 -88 -1849 88
rect -1895 -100 -1849 -88
rect -1799 88 -1753 100
rect -1799 -88 -1793 88
rect -1759 -88 -1753 88
rect -1799 -100 -1753 -88
rect -1703 88 -1657 100
rect -1703 -88 -1697 88
rect -1663 -88 -1657 88
rect -1703 -100 -1657 -88
rect -1607 88 -1561 100
rect -1607 -88 -1601 88
rect -1567 -88 -1561 88
rect -1607 -100 -1561 -88
rect -1511 88 -1465 100
rect -1511 -88 -1505 88
rect -1471 -88 -1465 88
rect -1511 -100 -1465 -88
rect -1415 88 -1369 100
rect -1415 -88 -1409 88
rect -1375 -88 -1369 88
rect -1415 -100 -1369 -88
rect -1319 88 -1273 100
rect -1319 -88 -1313 88
rect -1279 -88 -1273 88
rect -1319 -100 -1273 -88
rect -1223 88 -1177 100
rect -1223 -88 -1217 88
rect -1183 -88 -1177 88
rect -1223 -100 -1177 -88
rect -1127 88 -1081 100
rect -1127 -88 -1121 88
rect -1087 -88 -1081 88
rect -1127 -100 -1081 -88
rect -1031 88 -985 100
rect -1031 -88 -1025 88
rect -991 -88 -985 88
rect -1031 -100 -985 -88
rect -935 88 -889 100
rect -935 -88 -929 88
rect -895 -88 -889 88
rect -935 -100 -889 -88
rect -839 88 -793 100
rect -839 -88 -833 88
rect -799 -88 -793 88
rect -839 -100 -793 -88
rect -743 88 -697 100
rect -743 -88 -737 88
rect -703 -88 -697 88
rect -743 -100 -697 -88
rect -647 88 -601 100
rect -647 -88 -641 88
rect -607 -88 -601 88
rect -647 -100 -601 -88
rect -551 88 -505 100
rect -551 -88 -545 88
rect -511 -88 -505 88
rect -551 -100 -505 -88
rect -455 88 -409 100
rect -455 -88 -449 88
rect -415 -88 -409 88
rect -455 -100 -409 -88
rect -359 88 -313 100
rect -359 -88 -353 88
rect -319 -88 -313 88
rect -359 -100 -313 -88
rect -263 88 -217 100
rect -263 -88 -257 88
rect -223 -88 -217 88
rect -263 -100 -217 -88
rect -167 88 -121 100
rect -167 -88 -161 88
rect -127 -88 -121 88
rect -167 -100 -121 -88
rect -71 88 -25 100
rect -71 -88 -65 88
rect -31 -88 -25 88
rect -71 -100 -25 -88
rect 25 88 71 100
rect 25 -88 31 88
rect 65 -88 71 88
rect 25 -100 71 -88
rect 121 88 167 100
rect 121 -88 127 88
rect 161 -88 167 88
rect 121 -100 167 -88
rect 217 88 263 100
rect 217 -88 223 88
rect 257 -88 263 88
rect 217 -100 263 -88
rect 313 88 359 100
rect 313 -88 319 88
rect 353 -88 359 88
rect 313 -100 359 -88
rect 409 88 455 100
rect 409 -88 415 88
rect 449 -88 455 88
rect 409 -100 455 -88
rect 505 88 551 100
rect 505 -88 511 88
rect 545 -88 551 88
rect 505 -100 551 -88
rect 601 88 647 100
rect 601 -88 607 88
rect 641 -88 647 88
rect 601 -100 647 -88
rect 697 88 743 100
rect 697 -88 703 88
rect 737 -88 743 88
rect 697 -100 743 -88
rect 793 88 839 100
rect 793 -88 799 88
rect 833 -88 839 88
rect 793 -100 839 -88
rect 889 88 935 100
rect 889 -88 895 88
rect 929 -88 935 88
rect 889 -100 935 -88
rect 985 88 1031 100
rect 985 -88 991 88
rect 1025 -88 1031 88
rect 985 -100 1031 -88
rect 1081 88 1127 100
rect 1081 -88 1087 88
rect 1121 -88 1127 88
rect 1081 -100 1127 -88
rect 1177 88 1223 100
rect 1177 -88 1183 88
rect 1217 -88 1223 88
rect 1177 -100 1223 -88
rect 1273 88 1319 100
rect 1273 -88 1279 88
rect 1313 -88 1319 88
rect 1273 -100 1319 -88
rect 1369 88 1415 100
rect 1369 -88 1375 88
rect 1409 -88 1415 88
rect 1369 -100 1415 -88
rect 1465 88 1511 100
rect 1465 -88 1471 88
rect 1505 -88 1511 88
rect 1465 -100 1511 -88
rect 1561 88 1607 100
rect 1561 -88 1567 88
rect 1601 -88 1607 88
rect 1561 -100 1607 -88
rect 1657 88 1703 100
rect 1657 -88 1663 88
rect 1697 -88 1703 88
rect 1657 -100 1703 -88
rect 1753 88 1799 100
rect 1753 -88 1759 88
rect 1793 -88 1799 88
rect 1753 -100 1799 -88
rect 1849 88 1895 100
rect 1849 -88 1855 88
rect 1889 -88 1895 88
rect 1849 -100 1895 -88
rect 1945 88 1991 100
rect 1945 -88 1951 88
rect 1985 -88 1991 88
rect 1945 -100 1991 -88
rect 2041 88 2087 100
rect 2041 -88 2047 88
rect 2081 -88 2087 88
rect 2041 -100 2087 -88
rect 2137 88 2183 100
rect 2137 -88 2143 88
rect 2177 -88 2183 88
rect 2137 -100 2183 -88
rect 2233 88 2279 100
rect 2233 -88 2239 88
rect 2273 -88 2279 88
rect 2233 -100 2279 -88
rect 2329 88 2375 100
rect 2329 -88 2335 88
rect 2369 -88 2375 88
rect 2329 -100 2375 -88
rect 2425 88 2471 100
rect 2425 -88 2431 88
rect 2465 -88 2471 88
rect 2425 -100 2471 -88
rect 2521 88 2567 100
rect 2521 -88 2527 88
rect 2561 -88 2567 88
rect 2521 -100 2567 -88
rect 2617 88 2663 100
rect 2617 -88 2623 88
rect 2657 -88 2663 88
rect 2617 -100 2663 -88
rect 2713 88 2759 100
rect 2713 -88 2719 88
rect 2753 -88 2759 88
rect 2713 -100 2759 -88
rect 2809 88 2855 100
rect 2809 -88 2815 88
rect 2849 -88 2855 88
rect 2809 -100 2855 -88
rect 2905 88 2951 100
rect 2905 -88 2911 88
rect 2945 -88 2951 88
rect 2905 -100 2951 -88
rect -2909 -138 -2851 -132
rect -2909 -172 -2897 -138
rect -2863 -172 -2851 -138
rect -2909 -178 -2851 -172
rect -2717 -138 -2659 -132
rect -2717 -172 -2705 -138
rect -2671 -172 -2659 -138
rect -2717 -178 -2659 -172
rect -2525 -138 -2467 -132
rect -2525 -172 -2513 -138
rect -2479 -172 -2467 -138
rect -2525 -178 -2467 -172
rect -2333 -138 -2275 -132
rect -2333 -172 -2321 -138
rect -2287 -172 -2275 -138
rect -2333 -178 -2275 -172
rect -2141 -138 -2083 -132
rect -2141 -172 -2129 -138
rect -2095 -172 -2083 -138
rect -2141 -178 -2083 -172
rect -1949 -138 -1891 -132
rect -1949 -172 -1937 -138
rect -1903 -172 -1891 -138
rect -1949 -178 -1891 -172
rect -1757 -138 -1699 -132
rect -1757 -172 -1745 -138
rect -1711 -172 -1699 -138
rect -1757 -178 -1699 -172
rect -1565 -138 -1507 -132
rect -1565 -172 -1553 -138
rect -1519 -172 -1507 -138
rect -1565 -178 -1507 -172
rect -1373 -138 -1315 -132
rect -1373 -172 -1361 -138
rect -1327 -172 -1315 -138
rect -1373 -178 -1315 -172
rect -1181 -138 -1123 -132
rect -1181 -172 -1169 -138
rect -1135 -172 -1123 -138
rect -1181 -178 -1123 -172
rect -989 -138 -931 -132
rect -989 -172 -977 -138
rect -943 -172 -931 -138
rect -989 -178 -931 -172
rect -797 -138 -739 -132
rect -797 -172 -785 -138
rect -751 -172 -739 -138
rect -797 -178 -739 -172
rect -605 -138 -547 -132
rect -605 -172 -593 -138
rect -559 -172 -547 -138
rect -605 -178 -547 -172
rect -413 -138 -355 -132
rect -413 -172 -401 -138
rect -367 -172 -355 -138
rect -413 -178 -355 -172
rect -221 -138 -163 -132
rect -221 -172 -209 -138
rect -175 -172 -163 -138
rect -221 -178 -163 -172
rect -29 -138 29 -132
rect -29 -172 -17 -138
rect 17 -172 29 -138
rect -29 -178 29 -172
rect 163 -138 221 -132
rect 163 -172 175 -138
rect 209 -172 221 -138
rect 163 -178 221 -172
rect 355 -138 413 -132
rect 355 -172 367 -138
rect 401 -172 413 -138
rect 355 -178 413 -172
rect 547 -138 605 -132
rect 547 -172 559 -138
rect 593 -172 605 -138
rect 547 -178 605 -172
rect 739 -138 797 -132
rect 739 -172 751 -138
rect 785 -172 797 -138
rect 739 -178 797 -172
rect 931 -138 989 -132
rect 931 -172 943 -138
rect 977 -172 989 -138
rect 931 -178 989 -172
rect 1123 -138 1181 -132
rect 1123 -172 1135 -138
rect 1169 -172 1181 -138
rect 1123 -178 1181 -172
rect 1315 -138 1373 -132
rect 1315 -172 1327 -138
rect 1361 -172 1373 -138
rect 1315 -178 1373 -172
rect 1507 -138 1565 -132
rect 1507 -172 1519 -138
rect 1553 -172 1565 -138
rect 1507 -178 1565 -172
rect 1699 -138 1757 -132
rect 1699 -172 1711 -138
rect 1745 -172 1757 -138
rect 1699 -178 1757 -172
rect 1891 -138 1949 -132
rect 1891 -172 1903 -138
rect 1937 -172 1949 -138
rect 1891 -178 1949 -172
rect 2083 -138 2141 -132
rect 2083 -172 2095 -138
rect 2129 -172 2141 -138
rect 2083 -178 2141 -172
rect 2275 -138 2333 -132
rect 2275 -172 2287 -138
rect 2321 -172 2333 -138
rect 2275 -178 2333 -172
rect 2467 -138 2525 -132
rect 2467 -172 2479 -138
rect 2513 -172 2525 -138
rect 2467 -178 2525 -172
rect 2659 -138 2717 -132
rect 2659 -172 2671 -138
rect 2705 -172 2717 -138
rect 2659 -178 2717 -172
rect 2851 -138 2909 -132
rect 2851 -172 2863 -138
rect 2897 -172 2909 -138
rect 2851 -178 2909 -172
<< properties >>
string gencell sky130_fd_pr__nfet_01v8_lvt
string library sky130
string parameters w 1.0 l 0.15 m 1 nf 61 diffcov 100 polycov 100 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
