magic
tech sky130A
magscale 1 2
timestamp 1671746299
<< metal3 >>
rect -450 -500 449 500
<< mimcap >>
rect -350 360 250 400
rect -350 -360 -310 360
rect 210 -360 250 360
rect -350 -400 250 -360
<< mimcapcontact >>
rect -310 -360 210 360
<< metal4 >>
rect -311 360 211 361
rect -311 -360 -310 360
rect 210 -360 211 360
rect -311 -361 211 -360
<< properties >>
string FIXED_BBOX -450 -500 350 500
string gencell sky130_fd_pr__cap_mim_m3_1
string library sky130
string parameters w 3.0 l 4.0 val 26.66 carea 2.00 cperi 0.19 nx 1 ny 1 dummy 0 square 0 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 1 tconnect 1 ccov 100
<< end >>
