magic
tech sky130A
magscale 1 2
timestamp 1672092821
<< nwell >>
rect -1768 -538 1766 536
<< pmoslvt >>
rect -1572 117 -1502 317
rect -1444 117 -1374 317
rect -1316 117 -1246 317
rect -1188 117 -1118 317
rect -1060 117 -990 317
rect -932 117 -862 317
rect -804 117 -734 317
rect -676 117 -606 317
rect -548 117 -478 317
rect -420 117 -350 317
rect -292 117 -222 317
rect -164 117 -94 317
rect -36 117 34 317
rect 92 117 162 317
rect 220 117 290 317
rect 348 117 418 317
rect 476 117 546 317
rect 604 117 674 317
rect 732 117 802 317
rect 860 117 930 317
rect 988 117 1058 317
rect 1116 117 1186 317
rect 1244 117 1314 317
rect 1372 117 1442 317
rect 1500 117 1570 317
rect -1572 -319 -1502 -119
rect -1444 -319 -1374 -119
rect -1316 -319 -1246 -119
rect -1188 -319 -1118 -119
rect -1060 -319 -990 -119
rect -932 -319 -862 -119
rect -804 -319 -734 -119
rect -676 -319 -606 -119
rect -548 -319 -478 -119
rect -420 -319 -350 -119
rect -292 -319 -222 -119
rect -164 -319 -94 -119
rect -36 -319 34 -119
rect 92 -319 162 -119
rect 220 -319 290 -119
rect 348 -319 418 -119
rect 476 -319 546 -119
rect 604 -319 674 -119
rect 732 -319 802 -119
rect 860 -319 930 -119
rect 988 -319 1058 -119
rect 1116 -319 1186 -119
rect 1244 -319 1314 -119
rect 1372 -319 1442 -119
rect 1500 -319 1570 -119
<< pdiff >>
rect -1630 305 -1572 317
rect -1630 129 -1618 305
rect -1584 129 -1572 305
rect -1630 117 -1572 129
rect -1502 305 -1444 317
rect -1502 129 -1490 305
rect -1456 129 -1444 305
rect -1502 117 -1444 129
rect -1374 305 -1316 317
rect -1374 129 -1362 305
rect -1328 129 -1316 305
rect -1374 117 -1316 129
rect -1246 305 -1188 317
rect -1246 129 -1234 305
rect -1200 129 -1188 305
rect -1246 117 -1188 129
rect -1118 305 -1060 317
rect -1118 129 -1106 305
rect -1072 129 -1060 305
rect -1118 117 -1060 129
rect -990 305 -932 317
rect -990 129 -978 305
rect -944 129 -932 305
rect -990 117 -932 129
rect -862 305 -804 317
rect -862 129 -850 305
rect -816 129 -804 305
rect -862 117 -804 129
rect -734 305 -676 317
rect -734 129 -722 305
rect -688 129 -676 305
rect -734 117 -676 129
rect -606 305 -548 317
rect -606 129 -594 305
rect -560 129 -548 305
rect -606 117 -548 129
rect -478 305 -420 317
rect -478 129 -466 305
rect -432 129 -420 305
rect -478 117 -420 129
rect -350 305 -292 317
rect -350 129 -338 305
rect -304 129 -292 305
rect -350 117 -292 129
rect -222 305 -164 317
rect -222 129 -210 305
rect -176 129 -164 305
rect -222 117 -164 129
rect -94 305 -36 317
rect -94 129 -82 305
rect -48 129 -36 305
rect -94 117 -36 129
rect 34 305 92 317
rect 34 129 46 305
rect 80 129 92 305
rect 34 117 92 129
rect 162 305 220 317
rect 162 129 174 305
rect 208 129 220 305
rect 162 117 220 129
rect 290 305 348 317
rect 290 129 302 305
rect 336 129 348 305
rect 290 117 348 129
rect 418 305 476 317
rect 418 129 430 305
rect 464 129 476 305
rect 418 117 476 129
rect 546 305 604 317
rect 546 129 558 305
rect 592 129 604 305
rect 546 117 604 129
rect 674 305 732 317
rect 674 129 686 305
rect 720 129 732 305
rect 674 117 732 129
rect 802 305 860 317
rect 802 129 814 305
rect 848 129 860 305
rect 802 117 860 129
rect 930 305 988 317
rect 930 129 942 305
rect 976 129 988 305
rect 930 117 988 129
rect 1058 305 1116 317
rect 1058 129 1070 305
rect 1104 129 1116 305
rect 1058 117 1116 129
rect 1186 305 1244 317
rect 1186 129 1198 305
rect 1232 129 1244 305
rect 1186 117 1244 129
rect 1314 305 1372 317
rect 1314 129 1326 305
rect 1360 129 1372 305
rect 1314 117 1372 129
rect 1442 305 1500 317
rect 1442 129 1454 305
rect 1488 129 1500 305
rect 1442 117 1500 129
rect 1570 305 1628 317
rect 1570 129 1582 305
rect 1616 129 1628 305
rect 1570 117 1628 129
rect -1630 -131 -1572 -119
rect -1630 -307 -1618 -131
rect -1584 -307 -1572 -131
rect -1630 -319 -1572 -307
rect -1502 -131 -1444 -119
rect -1502 -307 -1490 -131
rect -1456 -307 -1444 -131
rect -1502 -319 -1444 -307
rect -1374 -131 -1316 -119
rect -1374 -307 -1362 -131
rect -1328 -307 -1316 -131
rect -1374 -319 -1316 -307
rect -1246 -131 -1188 -119
rect -1246 -307 -1234 -131
rect -1200 -307 -1188 -131
rect -1246 -319 -1188 -307
rect -1118 -131 -1060 -119
rect -1118 -307 -1106 -131
rect -1072 -307 -1060 -131
rect -1118 -319 -1060 -307
rect -990 -131 -932 -119
rect -990 -307 -978 -131
rect -944 -307 -932 -131
rect -990 -319 -932 -307
rect -862 -131 -804 -119
rect -862 -307 -850 -131
rect -816 -307 -804 -131
rect -862 -319 -804 -307
rect -734 -131 -676 -119
rect -734 -307 -722 -131
rect -688 -307 -676 -131
rect -734 -319 -676 -307
rect -606 -131 -548 -119
rect -606 -307 -594 -131
rect -560 -307 -548 -131
rect -606 -319 -548 -307
rect -478 -131 -420 -119
rect -478 -307 -466 -131
rect -432 -307 -420 -131
rect -478 -319 -420 -307
rect -350 -131 -292 -119
rect -350 -307 -338 -131
rect -304 -307 -292 -131
rect -350 -319 -292 -307
rect -222 -131 -164 -119
rect -222 -307 -210 -131
rect -176 -307 -164 -131
rect -222 -319 -164 -307
rect -94 -131 -36 -119
rect -94 -307 -82 -131
rect -48 -307 -36 -131
rect -94 -319 -36 -307
rect 34 -131 92 -119
rect 34 -307 46 -131
rect 80 -307 92 -131
rect 34 -319 92 -307
rect 162 -131 220 -119
rect 162 -307 174 -131
rect 208 -307 220 -131
rect 162 -319 220 -307
rect 290 -131 348 -119
rect 290 -307 302 -131
rect 336 -307 348 -131
rect 290 -319 348 -307
rect 418 -131 476 -119
rect 418 -307 430 -131
rect 464 -307 476 -131
rect 418 -319 476 -307
rect 546 -131 604 -119
rect 546 -307 558 -131
rect 592 -307 604 -131
rect 546 -319 604 -307
rect 674 -131 732 -119
rect 674 -307 686 -131
rect 720 -307 732 -131
rect 674 -319 732 -307
rect 802 -131 860 -119
rect 802 -307 814 -131
rect 848 -307 860 -131
rect 802 -319 860 -307
rect 930 -131 988 -119
rect 930 -307 942 -131
rect 976 -307 988 -131
rect 930 -319 988 -307
rect 1058 -131 1116 -119
rect 1058 -307 1070 -131
rect 1104 -307 1116 -131
rect 1058 -319 1116 -307
rect 1186 -131 1244 -119
rect 1186 -307 1198 -131
rect 1232 -307 1244 -131
rect 1186 -319 1244 -307
rect 1314 -131 1372 -119
rect 1314 -307 1326 -131
rect 1360 -307 1372 -131
rect 1314 -319 1372 -307
rect 1442 -131 1500 -119
rect 1442 -307 1454 -131
rect 1488 -307 1500 -131
rect 1442 -319 1500 -307
rect 1570 -131 1628 -119
rect 1570 -307 1582 -131
rect 1616 -307 1628 -131
rect 1570 -319 1628 -307
<< pdiffc >>
rect -1618 129 -1584 305
rect -1490 129 -1456 305
rect -1362 129 -1328 305
rect -1234 129 -1200 305
rect -1106 129 -1072 305
rect -978 129 -944 305
rect -850 129 -816 305
rect -722 129 -688 305
rect -594 129 -560 305
rect -466 129 -432 305
rect -338 129 -304 305
rect -210 129 -176 305
rect -82 129 -48 305
rect 46 129 80 305
rect 174 129 208 305
rect 302 129 336 305
rect 430 129 464 305
rect 558 129 592 305
rect 686 129 720 305
rect 814 129 848 305
rect 942 129 976 305
rect 1070 129 1104 305
rect 1198 129 1232 305
rect 1326 129 1360 305
rect 1454 129 1488 305
rect 1582 129 1616 305
rect -1618 -307 -1584 -131
rect -1490 -307 -1456 -131
rect -1362 -307 -1328 -131
rect -1234 -307 -1200 -131
rect -1106 -307 -1072 -131
rect -978 -307 -944 -131
rect -850 -307 -816 -131
rect -722 -307 -688 -131
rect -594 -307 -560 -131
rect -466 -307 -432 -131
rect -338 -307 -304 -131
rect -210 -307 -176 -131
rect -82 -307 -48 -131
rect 46 -307 80 -131
rect 174 -307 208 -131
rect 302 -307 336 -131
rect 430 -307 464 -131
rect 558 -307 592 -131
rect 686 -307 720 -131
rect 814 -307 848 -131
rect 942 -307 976 -131
rect 1070 -307 1104 -131
rect 1198 -307 1232 -131
rect 1326 -307 1360 -131
rect 1454 -307 1488 -131
rect 1582 -307 1616 -131
<< nsubdiff >>
rect -1732 466 -1636 500
rect 1634 466 1730 500
rect -1732 404 -1698 466
rect 1696 404 1730 466
rect -1732 -468 -1698 -406
rect 1696 -468 1730 -406
rect -1732 -502 -1636 -468
rect 1634 -502 1730 -468
<< nsubdiffcont >>
rect -1636 466 1634 500
rect -1732 -406 -1698 404
rect 1696 -406 1730 404
rect -1636 -502 1634 -468
<< poly >>
rect -1572 317 -1502 414
rect -1444 317 -1374 414
rect -1316 317 -1246 414
rect -1188 317 -1118 414
rect -1060 317 -990 414
rect -932 317 -862 414
rect -804 317 -734 414
rect -676 317 -606 414
rect -548 317 -478 414
rect -420 317 -350 414
rect -292 317 -222 414
rect -164 317 -94 414
rect -36 317 34 414
rect 92 317 162 414
rect 220 317 290 414
rect 348 317 418 414
rect 476 317 546 414
rect 604 317 674 414
rect 732 317 802 414
rect 860 317 930 414
rect 988 317 1058 414
rect 1116 317 1186 414
rect 1244 317 1314 414
rect 1372 317 1442 414
rect 1500 317 1570 414
rect -1572 -119 -1502 117
rect -1444 -119 -1374 117
rect -1316 -119 -1246 117
rect -1188 -119 -1118 117
rect -1060 -119 -990 117
rect -932 -119 -862 117
rect -804 -119 -734 117
rect -676 -119 -606 117
rect -548 -119 -478 117
rect -420 -119 -350 117
rect -292 -119 -222 117
rect -164 -119 -94 117
rect -36 -119 34 117
rect 92 -119 162 117
rect 220 -119 290 117
rect 348 -119 418 117
rect 476 -119 546 117
rect 604 -119 674 117
rect 732 -119 802 117
rect 860 -119 930 117
rect 988 -119 1058 117
rect 1116 -119 1186 117
rect 1244 -119 1314 117
rect 1372 -119 1442 117
rect 1500 -119 1570 117
rect -1572 -356 -1502 -319
rect -1444 -356 -1374 -319
rect -1316 -356 -1246 -319
rect -1188 -356 -1118 -319
rect -1060 -356 -990 -319
rect -932 -356 -862 -319
rect -804 -356 -734 -319
rect -676 -356 -606 -319
rect -548 -356 -478 -319
rect -420 -356 -350 -319
rect -292 -356 -222 -319
rect -164 -356 -94 -319
rect -36 -356 34 -319
rect 92 -356 162 -319
rect 220 -356 290 -319
rect 348 -356 418 -319
rect 476 -356 546 -319
rect 604 -356 674 -319
rect 732 -356 802 -319
rect 860 -356 930 -319
rect 988 -356 1058 -319
rect 1116 -356 1186 -319
rect 1244 -356 1314 -319
rect 1372 -356 1442 -319
rect 1500 -356 1570 -319
rect -1680 -374 1570 -356
rect -1680 -408 -1644 -374
rect -1596 -408 1570 -374
rect -1680 -432 1570 -408
<< polycont >>
rect -1644 -408 -1596 -374
<< locali >>
rect -1732 466 -1636 500
rect 1634 466 1730 500
rect -1732 404 -1698 466
rect 1696 404 1730 466
rect -1618 305 -1584 321
rect -1618 113 -1584 129
rect -1490 305 -1456 321
rect -1490 113 -1456 129
rect -1362 305 -1328 321
rect -1362 113 -1328 129
rect -1234 305 -1200 321
rect -1234 113 -1200 129
rect -1106 305 -1072 321
rect -1106 113 -1072 129
rect -978 305 -944 321
rect -978 113 -944 129
rect -850 305 -816 321
rect -850 113 -816 129
rect -722 305 -688 321
rect -722 113 -688 129
rect -594 305 -560 321
rect -594 113 -560 129
rect -466 305 -432 321
rect -466 113 -432 129
rect -338 305 -304 321
rect -338 113 -304 129
rect -210 305 -176 321
rect -210 113 -176 129
rect -82 305 -48 321
rect -82 113 -48 129
rect 46 305 80 321
rect 46 113 80 129
rect 174 305 208 321
rect 174 113 208 129
rect 302 305 336 321
rect 302 113 336 129
rect 430 305 464 321
rect 430 113 464 129
rect 558 305 592 321
rect 558 113 592 129
rect 686 305 720 321
rect 686 113 720 129
rect 814 305 848 321
rect 814 113 848 129
rect 942 305 976 321
rect 942 113 976 129
rect 1070 305 1104 321
rect 1070 113 1104 129
rect 1198 305 1232 321
rect 1198 113 1232 129
rect 1326 305 1360 321
rect 1326 113 1360 129
rect 1454 305 1488 321
rect 1454 113 1488 129
rect 1582 305 1616 321
rect 1582 113 1616 129
rect -1618 -131 -1584 -115
rect -1618 -323 -1584 -307
rect -1490 -131 -1456 -115
rect -1490 -323 -1456 -307
rect -1362 -131 -1328 -115
rect -1362 -323 -1328 -307
rect -1234 -131 -1200 -115
rect -1234 -323 -1200 -307
rect -1106 -131 -1072 -115
rect -1106 -323 -1072 -307
rect -978 -131 -944 -115
rect -978 -323 -944 -307
rect -850 -131 -816 -115
rect -850 -323 -816 -307
rect -722 -131 -688 -115
rect -722 -323 -688 -307
rect -594 -131 -560 -115
rect -594 -323 -560 -307
rect -466 -131 -432 -115
rect -466 -323 -432 -307
rect -338 -131 -304 -115
rect -338 -323 -304 -307
rect -210 -131 -176 -115
rect -210 -323 -176 -307
rect -82 -131 -48 -115
rect -82 -323 -48 -307
rect 46 -131 80 -115
rect 46 -323 80 -307
rect 174 -131 208 -115
rect 174 -323 208 -307
rect 302 -131 336 -115
rect 302 -323 336 -307
rect 430 -131 464 -115
rect 430 -323 464 -307
rect 558 -131 592 -115
rect 558 -323 592 -307
rect 686 -131 720 -115
rect 686 -323 720 -307
rect 814 -131 848 -115
rect 814 -323 848 -307
rect 942 -131 976 -115
rect 942 -323 976 -307
rect 1070 -131 1104 -115
rect 1070 -323 1104 -307
rect 1198 -131 1232 -115
rect 1198 -323 1232 -307
rect 1326 -131 1360 -115
rect 1326 -323 1360 -307
rect 1454 -131 1488 -115
rect 1454 -323 1488 -307
rect 1582 -131 1616 -115
rect 1582 -323 1616 -307
rect -1732 -468 -1698 -406
rect -1660 -368 -1580 -360
rect -1660 -416 -1652 -368
rect -1588 -416 -1580 -368
rect -1660 -424 -1580 -416
rect 1696 -468 1730 -406
rect -1732 -502 -1636 -468
rect 1634 -502 1730 -468
<< viali >>
rect -1618 129 -1584 305
rect -1490 129 -1456 305
rect -1362 129 -1328 305
rect -1234 129 -1200 305
rect -1106 129 -1072 305
rect -978 129 -944 305
rect -850 129 -816 305
rect -722 129 -688 305
rect -594 129 -560 305
rect -466 129 -432 305
rect -338 129 -304 305
rect -210 129 -176 305
rect -82 129 -48 305
rect 46 129 80 305
rect 174 129 208 305
rect 302 129 336 305
rect 430 129 464 305
rect 558 129 592 305
rect 686 129 720 305
rect 814 129 848 305
rect 942 129 976 305
rect 1070 129 1104 305
rect 1198 129 1232 305
rect 1326 129 1360 305
rect 1454 129 1488 305
rect 1582 129 1616 305
rect -1618 -307 -1584 -131
rect -1490 -307 -1456 -131
rect -1362 -307 -1328 -131
rect -1234 -307 -1200 -131
rect -1106 -307 -1072 -131
rect -978 -307 -944 -131
rect -850 -307 -816 -131
rect -722 -307 -688 -131
rect -594 -307 -560 -131
rect -466 -307 -432 -131
rect -338 -307 -304 -131
rect -210 -307 -176 -131
rect -82 -307 -48 -131
rect 46 -307 80 -131
rect 174 -307 208 -131
rect 302 -307 336 -131
rect 430 -307 464 -131
rect 558 -307 592 -131
rect 686 -307 720 -131
rect 814 -307 848 -131
rect 942 -307 976 -131
rect 1070 -307 1104 -131
rect 1198 -307 1232 -131
rect 1326 -307 1360 -131
rect 1454 -307 1488 -131
rect 1582 -307 1616 -131
rect -1652 -374 -1588 -368
rect -1652 -408 -1644 -374
rect -1644 -408 -1596 -374
rect -1596 -408 -1588 -374
rect -1652 -416 -1588 -408
<< metal1 >>
rect -1630 444 -1572 456
rect -1630 336 -1628 444
rect -1574 336 -1572 444
rect -1630 314 -1572 336
rect -1374 444 -1316 456
rect -1374 336 -1372 444
rect -1318 336 -1316 444
rect -1624 305 -1578 314
rect -1624 129 -1618 305
rect -1584 129 -1578 305
rect -1624 -131 -1578 129
rect -1496 305 -1450 317
rect -1374 314 -1316 336
rect -1118 444 -1060 456
rect -1118 336 -1116 444
rect -1062 336 -1060 444
rect -1496 129 -1490 305
rect -1456 129 -1450 305
rect -1496 118 -1450 129
rect -1368 305 -1322 314
rect -1368 129 -1362 305
rect -1328 129 -1322 305
rect -1502 78 -1444 118
rect -1502 -80 -1498 78
rect -1446 -80 -1444 78
rect -1502 -120 -1444 -80
rect -1624 -307 -1618 -131
rect -1584 -307 -1578 -131
rect -1624 -319 -1578 -307
rect -1496 -131 -1450 -120
rect -1496 -307 -1490 -131
rect -1456 -307 -1450 -131
rect -1496 -319 -1450 -307
rect -1368 -131 -1322 129
rect -1240 305 -1194 317
rect -1118 314 -1060 336
rect -862 444 -804 456
rect -862 336 -860 444
rect -806 336 -804 444
rect -1240 129 -1234 305
rect -1200 129 -1194 305
rect -1240 118 -1194 129
rect -1112 305 -1066 314
rect -1112 129 -1106 305
rect -1072 129 -1066 305
rect -1246 78 -1188 118
rect -1246 -80 -1242 78
rect -1190 -80 -1188 78
rect -1246 -120 -1188 -80
rect -1368 -307 -1362 -131
rect -1328 -307 -1322 -131
rect -1368 -319 -1322 -307
rect -1240 -131 -1194 -120
rect -1240 -307 -1234 -131
rect -1200 -307 -1194 -131
rect -1240 -319 -1194 -307
rect -1112 -131 -1066 129
rect -984 305 -938 317
rect -862 314 -804 336
rect -606 444 -548 456
rect -606 336 -604 444
rect -550 336 -548 444
rect -984 129 -978 305
rect -944 129 -938 305
rect -984 118 -938 129
rect -856 305 -810 314
rect -856 129 -850 305
rect -816 129 -810 305
rect -990 78 -932 118
rect -990 -80 -986 78
rect -934 -80 -932 78
rect -990 -120 -932 -80
rect -1112 -307 -1106 -131
rect -1072 -307 -1066 -131
rect -1112 -319 -1066 -307
rect -984 -131 -938 -120
rect -984 -307 -978 -131
rect -944 -307 -938 -131
rect -984 -319 -938 -307
rect -856 -131 -810 129
rect -728 305 -682 317
rect -606 314 -548 336
rect -350 444 -292 456
rect -350 336 -348 444
rect -294 336 -292 444
rect -728 129 -722 305
rect -688 129 -682 305
rect -728 118 -682 129
rect -600 305 -554 314
rect -600 129 -594 305
rect -560 129 -554 305
rect -734 78 -676 118
rect -734 -80 -730 78
rect -678 -80 -676 78
rect -734 -120 -676 -80
rect -856 -307 -850 -131
rect -816 -307 -810 -131
rect -856 -319 -810 -307
rect -728 -131 -682 -120
rect -728 -307 -722 -131
rect -688 -307 -682 -131
rect -728 -319 -682 -307
rect -600 -131 -554 129
rect -472 305 -426 317
rect -350 314 -292 336
rect -94 444 -36 456
rect -94 336 -92 444
rect -38 336 -36 444
rect -472 129 -466 305
rect -432 129 -426 305
rect -472 118 -426 129
rect -344 305 -298 314
rect -344 129 -338 305
rect -304 129 -298 305
rect -478 78 -420 118
rect -478 -80 -474 78
rect -422 -80 -420 78
rect -478 -120 -420 -80
rect -600 -307 -594 -131
rect -560 -307 -554 -131
rect -600 -319 -554 -307
rect -472 -131 -426 -120
rect -472 -307 -466 -131
rect -432 -307 -426 -131
rect -472 -319 -426 -307
rect -344 -131 -298 129
rect -216 305 -170 317
rect -94 314 -36 336
rect 162 444 220 456
rect 162 336 164 444
rect 218 336 220 444
rect -216 129 -210 305
rect -176 129 -170 305
rect -216 118 -170 129
rect -88 305 -42 314
rect -88 129 -82 305
rect -48 129 -42 305
rect -222 78 -164 118
rect -222 -80 -218 78
rect -166 -80 -164 78
rect -222 -120 -164 -80
rect -344 -307 -338 -131
rect -304 -307 -298 -131
rect -344 -319 -298 -307
rect -216 -131 -170 -120
rect -216 -307 -210 -131
rect -176 -307 -170 -131
rect -216 -319 -170 -307
rect -88 -131 -42 129
rect 40 305 86 317
rect 162 314 220 336
rect 418 444 476 456
rect 418 336 420 444
rect 474 336 476 444
rect 40 129 46 305
rect 80 129 86 305
rect 40 118 86 129
rect 168 305 214 314
rect 168 129 174 305
rect 208 129 214 305
rect 34 78 92 118
rect 34 -80 38 78
rect 90 -80 92 78
rect 34 -120 92 -80
rect -88 -307 -82 -131
rect -48 -307 -42 -131
rect -88 -319 -42 -307
rect 40 -131 86 -120
rect 40 -307 46 -131
rect 80 -307 86 -131
rect 40 -319 86 -307
rect 168 -131 214 129
rect 296 305 342 317
rect 418 314 476 336
rect 674 444 732 456
rect 674 336 676 444
rect 730 336 732 444
rect 296 129 302 305
rect 336 129 342 305
rect 296 118 342 129
rect 424 305 470 314
rect 424 129 430 305
rect 464 129 470 305
rect 290 78 348 118
rect 290 -80 294 78
rect 346 -80 348 78
rect 290 -120 348 -80
rect 168 -307 174 -131
rect 208 -307 214 -131
rect 168 -319 214 -307
rect 296 -131 342 -120
rect 296 -307 302 -131
rect 336 -307 342 -131
rect 296 -319 342 -307
rect 424 -131 470 129
rect 552 305 598 317
rect 674 314 732 336
rect 930 444 988 456
rect 930 336 932 444
rect 986 336 988 444
rect 552 129 558 305
rect 592 129 598 305
rect 552 118 598 129
rect 680 305 726 314
rect 680 129 686 305
rect 720 129 726 305
rect 546 78 604 118
rect 546 -80 550 78
rect 602 -80 604 78
rect 546 -120 604 -80
rect 424 -307 430 -131
rect 464 -307 470 -131
rect 424 -319 470 -307
rect 552 -131 598 -120
rect 552 -307 558 -131
rect 592 -307 598 -131
rect 552 -319 598 -307
rect 680 -131 726 129
rect 808 305 854 317
rect 930 314 988 336
rect 1186 444 1244 456
rect 1186 336 1188 444
rect 1242 336 1244 444
rect 808 129 814 305
rect 848 129 854 305
rect 808 118 854 129
rect 936 305 982 314
rect 936 129 942 305
rect 976 129 982 305
rect 802 78 860 118
rect 802 -80 806 78
rect 858 -80 860 78
rect 802 -120 860 -80
rect 680 -307 686 -131
rect 720 -307 726 -131
rect 680 -319 726 -307
rect 808 -131 854 -120
rect 808 -307 814 -131
rect 848 -307 854 -131
rect 808 -319 854 -307
rect 936 -131 982 129
rect 1064 305 1110 317
rect 1186 314 1244 336
rect 1442 444 1500 456
rect 1442 336 1444 444
rect 1498 336 1500 444
rect 1064 129 1070 305
rect 1104 129 1110 305
rect 1064 118 1110 129
rect 1192 305 1238 314
rect 1192 129 1198 305
rect 1232 129 1238 305
rect 1058 78 1116 118
rect 1058 -80 1062 78
rect 1114 -80 1116 78
rect 1058 -120 1116 -80
rect 936 -307 942 -131
rect 976 -307 982 -131
rect 936 -319 982 -307
rect 1064 -131 1110 -120
rect 1064 -307 1070 -131
rect 1104 -307 1110 -131
rect 1064 -319 1110 -307
rect 1192 -131 1238 129
rect 1320 305 1366 317
rect 1442 314 1500 336
rect 1320 129 1326 305
rect 1360 129 1366 305
rect 1320 118 1366 129
rect 1448 305 1494 314
rect 1448 129 1454 305
rect 1488 129 1494 305
rect 1314 78 1372 118
rect 1314 -80 1318 78
rect 1370 -80 1372 78
rect 1314 -120 1372 -80
rect 1192 -307 1198 -131
rect 1232 -307 1238 -131
rect 1192 -319 1238 -307
rect 1320 -131 1366 -120
rect 1320 -307 1326 -131
rect 1360 -307 1366 -131
rect 1320 -319 1366 -307
rect 1448 -131 1494 129
rect 1576 305 1622 317
rect 1576 129 1582 305
rect 1616 129 1622 305
rect 1576 118 1622 129
rect 1570 78 1628 118
rect 1570 -80 1574 78
rect 1626 -80 1628 78
rect 1570 -120 1628 -80
rect 1448 -307 1454 -131
rect 1488 -307 1494 -131
rect 1448 -319 1494 -307
rect 1576 -131 1622 -120
rect 1576 -307 1582 -131
rect 1616 -307 1622 -131
rect 1576 -319 1622 -307
rect -1680 -368 -1576 -356
rect -1680 -416 -1652 -368
rect -1588 -416 -1576 -368
rect -1680 -432 -1576 -416
<< via1 >>
rect -1628 336 -1574 444
rect -1372 336 -1318 444
rect -1116 336 -1062 444
rect -1498 -80 -1446 78
rect -860 336 -806 444
rect -1242 -80 -1190 78
rect -604 336 -550 444
rect -986 -80 -934 78
rect -348 336 -294 444
rect -730 -80 -678 78
rect -92 336 -38 444
rect -474 -80 -422 78
rect 164 336 218 444
rect -218 -80 -166 78
rect 420 336 474 444
rect 38 -80 90 78
rect 676 336 730 444
rect 294 -80 346 78
rect 932 336 986 444
rect 550 -80 602 78
rect 1188 336 1242 444
rect 806 -80 858 78
rect 1444 336 1498 444
rect 1062 -80 1114 78
rect 1318 -80 1370 78
rect 1574 -80 1626 78
<< metal2 >>
rect -1630 444 1628 614
rect -1630 336 -1628 444
rect -1574 336 -1372 444
rect -1318 336 -1116 444
rect -1062 336 -860 444
rect -806 336 -604 444
rect -550 336 -348 444
rect -294 336 -92 444
rect -38 336 164 444
rect 218 336 420 444
rect 474 336 676 444
rect 730 336 932 444
rect 986 336 1188 444
rect 1242 336 1444 444
rect 1498 336 1628 444
rect -1630 294 1628 336
rect -1630 78 1628 156
rect -1630 -80 -1498 78
rect -1446 -80 -1242 78
rect -1190 -80 -986 78
rect -934 -80 -730 78
rect -678 -80 -474 78
rect -422 -80 -218 78
rect -166 -80 38 78
rect 90 -80 294 78
rect 346 -80 550 78
rect 602 -80 806 78
rect 858 -80 1062 78
rect 1114 -80 1318 78
rect 1370 -80 1574 78
rect 1626 -80 1628 78
rect -1630 -164 1628 -80
<< properties >>
string FIXED_BBOX -1714 -484 1714 484
string gencell sky130_fd_pr__pfet_01v8_lvt
string library sky130
string parameters w 1.0 l 0.35 m 2 nf 25 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.35 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
