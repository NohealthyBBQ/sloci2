magic
tech sky130A
magscale 1 2
timestamp 1662690363
<< error_p >>
rect -159 -111 -97 -105
rect -31 -111 31 -105
rect 97 -111 159 -105
rect -159 -145 -147 -111
rect -31 -145 -19 -111
rect 97 -145 109 -111
rect -159 -151 -97 -145
rect -31 -151 31 -145
rect 97 -151 159 -145
<< nwell >>
rect -359 -284 359 284
<< pmoslvt >>
rect -163 -64 -93 136
rect -35 -64 35 136
rect 93 -64 163 136
<< pdiff >>
rect -221 124 -163 136
rect -221 -52 -209 124
rect -175 -52 -163 124
rect -221 -64 -163 -52
rect -93 124 -35 136
rect -93 -52 -81 124
rect -47 -52 -35 124
rect -93 -64 -35 -52
rect 35 124 93 136
rect 35 -52 47 124
rect 81 -52 93 124
rect 35 -64 93 -52
rect 163 124 221 136
rect 163 -52 175 124
rect 209 -52 221 124
rect 163 -64 221 -52
<< pdiffc >>
rect -209 -52 -175 124
rect -81 -52 -47 124
rect 47 -52 81 124
rect 175 -52 209 124
<< nsubdiff >>
rect -323 214 -227 248
rect 227 214 323 248
rect -323 151 -289 214
rect 289 151 323 214
rect -323 -214 -289 -151
rect 289 -214 323 -151
rect -323 -248 -227 -214
rect 227 -248 323 -214
<< nsubdiffcont >>
rect -227 214 227 248
rect -323 -151 -289 151
rect 289 -151 323 151
rect -227 -248 227 -214
<< poly >>
rect -163 136 -93 162
rect -35 136 35 162
rect 93 136 163 162
rect -163 -111 -93 -64
rect -163 -145 -147 -111
rect -109 -145 -93 -111
rect -163 -161 -93 -145
rect -35 -111 35 -64
rect -35 -145 -19 -111
rect 19 -145 35 -111
rect -35 -161 35 -145
rect 93 -111 163 -64
rect 93 -145 109 -111
rect 147 -145 163 -111
rect 93 -161 163 -145
<< polycont >>
rect -147 -145 -109 -111
rect -19 -145 19 -111
rect 109 -145 147 -111
<< locali >>
rect -323 214 -227 248
rect 227 214 323 248
rect -323 151 -289 214
rect 289 151 323 214
rect -209 124 -175 140
rect -209 -68 -175 -52
rect -81 124 -47 140
rect -81 -68 -47 -52
rect 47 124 81 140
rect 47 -68 81 -52
rect 175 124 209 140
rect 175 -68 209 -52
rect -163 -145 -147 -111
rect -109 -145 -93 -111
rect -35 -145 -19 -111
rect 19 -145 35 -111
rect 93 -145 109 -111
rect 147 -145 163 -111
rect -323 -214 -289 -151
rect 289 -214 323 -151
rect -323 -248 -227 -214
rect 227 -248 323 -214
<< viali >>
rect -209 -52 -175 124
rect -81 -52 -47 124
rect 47 -52 81 124
rect 175 -52 209 124
rect -147 -145 -109 -111
rect -19 -145 19 -111
rect 109 -145 147 -111
<< metal1 >>
rect -215 124 -169 136
rect -215 -52 -209 124
rect -175 -52 -169 124
rect -215 -64 -169 -52
rect -87 124 -41 136
rect -87 -52 -81 124
rect -47 -52 -41 124
rect -87 -64 -41 -52
rect 41 124 87 136
rect 41 -52 47 124
rect 81 -52 87 124
rect 41 -64 87 -52
rect 169 124 215 136
rect 169 -52 175 124
rect 209 -52 215 124
rect 169 -64 215 -52
rect -159 -111 -97 -105
rect -159 -145 -147 -111
rect -109 -145 -97 -111
rect -159 -151 -97 -145
rect -31 -111 31 -105
rect -31 -145 -19 -111
rect 19 -145 31 -111
rect -31 -151 31 -145
rect 97 -111 159 -105
rect 97 -145 109 -111
rect 147 -145 159 -111
rect 97 -151 159 -145
<< properties >>
string FIXED_BBOX -306 -231 306 231
string gencell sky130_fd_pr__pfet_01v8_lvt
string library sky130
string parameters w 1 l 0.35 m 1 nf 3 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 0 botc 1 poverlap 0 doverlap 1 lmin 0.35 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
