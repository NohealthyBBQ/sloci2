magic
tech sky130A
magscale 1 2
timestamp 1662404926
<< metal3 >>
rect -2150 3072 2149 3100
rect -2150 -3072 2065 3072
rect 2129 -3072 2149 3072
rect -2150 -3100 2149 -3072
<< via3 >>
rect 2065 -3072 2129 3072
<< mimcap >>
rect -2050 2960 1950 3000
rect -2050 -2960 -2010 2960
rect 1910 -2960 1950 2960
rect -2050 -3000 1950 -2960
<< mimcapcontact >>
rect -2010 -2960 1910 2960
<< metal4 >>
rect 2049 3072 2145 3088
rect -2011 2960 1911 2961
rect -2011 -2960 -2010 2960
rect 1910 -2960 1911 2960
rect -2011 -2961 1911 -2960
rect 2049 -3072 2065 3072
rect 2129 -3072 2145 3072
rect 2049 -3088 2145 -3072
<< properties >>
string FIXED_BBOX -2150 -3100 2050 3100
string gencell sky130_fd_pr__cap_mim_m3_1
string library sky130
string parameters w 20.0 l 30.0 val 1.219k carea 2.00 cperi 0.19 nx 1 ny 1 dummy 0 square 0 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 1 tconnect 1 ccov 100
<< end >>
