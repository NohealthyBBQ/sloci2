magic
tech sky130A
magscale 1 2
timestamp 1671746188
<< metal3 >>
rect -1350 -1700 1349 1700
<< mimcap >>
rect -1250 1560 1150 1600
rect -1250 -1560 -1210 1560
rect 1110 -1560 1150 1560
rect -1250 -1600 1150 -1560
<< mimcapcontact >>
rect -1210 -1560 1110 1560
<< metal4 >>
rect -1211 1560 1111 1561
rect -1211 -1560 -1210 1560
rect 1110 -1560 1111 1560
rect -1211 -1561 1111 -1560
<< properties >>
string FIXED_BBOX -1350 -1700 1250 1700
string gencell sky130_fd_pr__cap_mim_m3_1
string library sky130
string parameters w 12.0 l 16.0 val 394.64 carea 2.00 cperi 0.19 nx 1 ny 1 dummy 0 square 0 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 1 tconnect 1 ccov 100
<< end >>
