magic
tech sky130A
magscale 1 2
timestamp 1662404926
<< error_p >>
rect -365 172 -307 178
rect -173 172 -115 178
rect 19 172 77 178
rect 211 172 269 178
rect 403 172 461 178
rect -365 138 -353 172
rect -173 138 -161 172
rect 19 138 31 172
rect 211 138 223 172
rect 403 138 415 172
rect -365 132 -307 138
rect -173 132 -115 138
rect 19 132 77 138
rect 211 132 269 138
rect 403 132 461 138
rect -461 -138 -403 -132
rect -269 -138 -211 -132
rect -77 -138 -19 -132
rect 115 -138 173 -132
rect 307 -138 365 -132
rect -461 -172 -449 -138
rect -269 -172 -257 -138
rect -77 -172 -65 -138
rect 115 -172 127 -138
rect 307 -172 319 -138
rect -461 -178 -403 -172
rect -269 -178 -211 -172
rect -77 -178 -19 -172
rect 115 -178 173 -172
rect 307 -178 365 -172
<< pwell >>
rect -647 -310 647 310
<< nmoslvt >>
rect -447 -100 -417 100
rect -351 -100 -321 100
rect -255 -100 -225 100
rect -159 -100 -129 100
rect -63 -100 -33 100
rect 33 -100 63 100
rect 129 -100 159 100
rect 225 -100 255 100
rect 321 -100 351 100
rect 417 -100 447 100
<< ndiff >>
rect -509 88 -447 100
rect -509 -88 -497 88
rect -463 -88 -447 88
rect -509 -100 -447 -88
rect -417 88 -351 100
rect -417 -88 -401 88
rect -367 -88 -351 88
rect -417 -100 -351 -88
rect -321 88 -255 100
rect -321 -88 -305 88
rect -271 -88 -255 88
rect -321 -100 -255 -88
rect -225 88 -159 100
rect -225 -88 -209 88
rect -175 -88 -159 88
rect -225 -100 -159 -88
rect -129 88 -63 100
rect -129 -88 -113 88
rect -79 -88 -63 88
rect -129 -100 -63 -88
rect -33 88 33 100
rect -33 -88 -17 88
rect 17 -88 33 88
rect -33 -100 33 -88
rect 63 88 129 100
rect 63 -88 79 88
rect 113 -88 129 88
rect 63 -100 129 -88
rect 159 88 225 100
rect 159 -88 175 88
rect 209 -88 225 88
rect 159 -100 225 -88
rect 255 88 321 100
rect 255 -88 271 88
rect 305 -88 321 88
rect 255 -100 321 -88
rect 351 88 417 100
rect 351 -88 367 88
rect 401 -88 417 88
rect 351 -100 417 -88
rect 447 88 509 100
rect 447 -88 463 88
rect 497 -88 509 88
rect 447 -100 509 -88
<< ndiffc >>
rect -497 -88 -463 88
rect -401 -88 -367 88
rect -305 -88 -271 88
rect -209 -88 -175 88
rect -113 -88 -79 88
rect -17 -88 17 88
rect 79 -88 113 88
rect 175 -88 209 88
rect 271 -88 305 88
rect 367 -88 401 88
rect 463 -88 497 88
<< psubdiff >>
rect -611 240 -515 274
rect 515 240 611 274
rect -611 178 -577 240
rect 577 178 611 240
rect -611 -240 -577 -178
rect 577 -240 611 -178
rect -611 -274 -515 -240
rect 515 -274 611 -240
<< psubdiffcont >>
rect -515 240 515 274
rect -611 -178 -577 178
rect 577 -178 611 178
rect -515 -274 515 -240
<< poly >>
rect -369 172 -303 188
rect -369 138 -353 172
rect -319 138 -303 172
rect -447 100 -417 126
rect -369 122 -303 138
rect -177 172 -111 188
rect -177 138 -161 172
rect -127 138 -111 172
rect -351 100 -321 122
rect -255 100 -225 126
rect -177 122 -111 138
rect 15 172 81 188
rect 15 138 31 172
rect 65 138 81 172
rect -159 100 -129 122
rect -63 100 -33 126
rect 15 122 81 138
rect 207 172 273 188
rect 207 138 223 172
rect 257 138 273 172
rect 33 100 63 122
rect 129 100 159 126
rect 207 122 273 138
rect 399 172 465 188
rect 399 138 415 172
rect 449 138 465 172
rect 225 100 255 122
rect 321 100 351 126
rect 399 122 465 138
rect 417 100 447 122
rect -447 -122 -417 -100
rect -465 -138 -399 -122
rect -351 -126 -321 -100
rect -255 -122 -225 -100
rect -465 -172 -449 -138
rect -415 -172 -399 -138
rect -465 -188 -399 -172
rect -273 -138 -207 -122
rect -159 -126 -129 -100
rect -63 -122 -33 -100
rect -273 -172 -257 -138
rect -223 -172 -207 -138
rect -273 -188 -207 -172
rect -81 -138 -15 -122
rect 33 -126 63 -100
rect 129 -122 159 -100
rect -81 -172 -65 -138
rect -31 -172 -15 -138
rect -81 -188 -15 -172
rect 111 -138 177 -122
rect 225 -126 255 -100
rect 321 -122 351 -100
rect 111 -172 127 -138
rect 161 -172 177 -138
rect 111 -188 177 -172
rect 303 -138 369 -122
rect 417 -126 447 -100
rect 303 -172 319 -138
rect 353 -172 369 -138
rect 303 -188 369 -172
<< polycont >>
rect -353 138 -319 172
rect -161 138 -127 172
rect 31 138 65 172
rect 223 138 257 172
rect 415 138 449 172
rect -449 -172 -415 -138
rect -257 -172 -223 -138
rect -65 -172 -31 -138
rect 127 -172 161 -138
rect 319 -172 353 -138
<< locali >>
rect -611 240 -515 274
rect 515 240 611 274
rect -611 178 -577 240
rect 577 178 611 240
rect -369 138 -353 172
rect -319 138 -303 172
rect -177 138 -161 172
rect -127 138 -111 172
rect 15 138 31 172
rect 65 138 81 172
rect 207 138 223 172
rect 257 138 273 172
rect 399 138 415 172
rect 449 138 465 172
rect -497 88 -463 104
rect -497 -104 -463 -88
rect -401 88 -367 104
rect -401 -104 -367 -88
rect -305 88 -271 104
rect -305 -104 -271 -88
rect -209 88 -175 104
rect -209 -104 -175 -88
rect -113 88 -79 104
rect -113 -104 -79 -88
rect -17 88 17 104
rect -17 -104 17 -88
rect 79 88 113 104
rect 79 -104 113 -88
rect 175 88 209 104
rect 175 -104 209 -88
rect 271 88 305 104
rect 271 -104 305 -88
rect 367 88 401 104
rect 367 -104 401 -88
rect 463 88 497 104
rect 463 -104 497 -88
rect -465 -172 -449 -138
rect -415 -172 -399 -138
rect -273 -172 -257 -138
rect -223 -172 -207 -138
rect -81 -172 -65 -138
rect -31 -172 -15 -138
rect 111 -172 127 -138
rect 161 -172 177 -138
rect 303 -172 319 -138
rect 353 -172 369 -138
rect -611 -240 -577 -178
rect 577 -240 611 -178
rect -611 -274 -515 -240
rect 515 -274 611 -240
<< viali >>
rect -353 138 -319 172
rect -161 138 -127 172
rect 31 138 65 172
rect 223 138 257 172
rect 415 138 449 172
rect -497 -88 -463 88
rect -401 -88 -367 88
rect -305 -88 -271 88
rect -209 -88 -175 88
rect -113 -88 -79 88
rect -17 -88 17 88
rect 79 -88 113 88
rect 175 -88 209 88
rect 271 -88 305 88
rect 367 -88 401 88
rect 463 -88 497 88
rect -449 -172 -415 -138
rect -257 -172 -223 -138
rect -65 -172 -31 -138
rect 127 -172 161 -138
rect 319 -172 353 -138
<< metal1 >>
rect -365 172 -307 178
rect -365 138 -353 172
rect -319 138 -307 172
rect -365 132 -307 138
rect -173 172 -115 178
rect -173 138 -161 172
rect -127 138 -115 172
rect -173 132 -115 138
rect 19 172 77 178
rect 19 138 31 172
rect 65 138 77 172
rect 19 132 77 138
rect 211 172 269 178
rect 211 138 223 172
rect 257 138 269 172
rect 211 132 269 138
rect 403 172 461 178
rect 403 138 415 172
rect 449 138 461 172
rect 403 132 461 138
rect -503 88 -457 100
rect -503 -88 -497 88
rect -463 -88 -457 88
rect -503 -100 -457 -88
rect -407 88 -361 100
rect -407 -88 -401 88
rect -367 -88 -361 88
rect -407 -100 -361 -88
rect -311 88 -265 100
rect -311 -88 -305 88
rect -271 -88 -265 88
rect -311 -100 -265 -88
rect -215 88 -169 100
rect -215 -88 -209 88
rect -175 -88 -169 88
rect -215 -100 -169 -88
rect -119 88 -73 100
rect -119 -88 -113 88
rect -79 -88 -73 88
rect -119 -100 -73 -88
rect -23 88 23 100
rect -23 -88 -17 88
rect 17 -88 23 88
rect -23 -100 23 -88
rect 73 88 119 100
rect 73 -88 79 88
rect 113 -88 119 88
rect 73 -100 119 -88
rect 169 88 215 100
rect 169 -88 175 88
rect 209 -88 215 88
rect 169 -100 215 -88
rect 265 88 311 100
rect 265 -88 271 88
rect 305 -88 311 88
rect 265 -100 311 -88
rect 361 88 407 100
rect 361 -88 367 88
rect 401 -88 407 88
rect 361 -100 407 -88
rect 457 88 503 100
rect 457 -88 463 88
rect 497 -88 503 88
rect 457 -100 503 -88
rect -461 -138 -403 -132
rect -461 -172 -449 -138
rect -415 -172 -403 -138
rect -461 -178 -403 -172
rect -269 -138 -211 -132
rect -269 -172 -257 -138
rect -223 -172 -211 -138
rect -269 -178 -211 -172
rect -77 -138 -19 -132
rect -77 -172 -65 -138
rect -31 -172 -19 -138
rect -77 -178 -19 -172
rect 115 -138 173 -132
rect 115 -172 127 -138
rect 161 -172 173 -138
rect 115 -178 173 -172
rect 307 -138 365 -132
rect 307 -172 319 -138
rect 353 -172 365 -138
rect 307 -178 365 -172
<< properties >>
string FIXED_BBOX -594 -257 594 257
string gencell sky130_fd_pr__nfet_01v8_lvt
string library sky130
string parameters w 1.0 l 0.15 m 1 nf 10 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
