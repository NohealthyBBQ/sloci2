magic
tech sky130A
magscale 1 2
timestamp 1662983156
<< pwell >>
rect 53403 -7310 53408 -7308
<< ndiff >>
rect 53403 -7310 53408 -7308
<< locali >>
rect 48302 -6398 48426 -6396
rect 48302 -6542 48820 -6398
rect 68132 -6416 68246 -6400
rect 67728 -6536 68246 -6416
rect 68132 -6542 68246 -6536
rect 49802 -7670 49900 -7624
<< viali >>
rect 48274 -7764 48446 -7706
rect 49940 -7756 66588 -7664
rect 68120 -7768 68292 -7710
<< metal1 >>
rect 48934 -5718 49008 -5432
rect 67544 -5802 67616 -5516
rect 47244 -7752 47254 -6678
rect 47614 -7752 47624 -6678
rect 48194 -7112 48556 -6644
rect 49426 -6924 49436 -6872
rect 49488 -6924 49498 -6872
rect 49432 -7112 49484 -6924
rect 48194 -7202 49484 -7112
rect 48194 -7240 48556 -7202
rect 48190 -7640 48556 -7240
rect 49538 -7692 49590 -7036
rect 49672 -7312 49724 -6302
rect 51874 -6610 51904 -6358
rect 64088 -6610 64118 -6352
rect 51874 -6640 57930 -6610
rect 51874 -6920 51904 -6640
rect 52038 -6741 52048 -6689
rect 52100 -6741 52110 -6689
rect 52228 -6740 52238 -6688
rect 52290 -6740 52300 -6688
rect 52420 -6739 52430 -6687
rect 52482 -6739 52492 -6687
rect 52611 -6739 52621 -6687
rect 52673 -6739 52683 -6687
rect 52805 -6739 52815 -6687
rect 52867 -6739 52877 -6687
rect 52995 -6740 53005 -6688
rect 53057 -6740 53067 -6688
rect 53189 -6739 53199 -6687
rect 53251 -6739 53261 -6687
rect 53381 -6739 53391 -6687
rect 53443 -6739 53453 -6687
rect 53572 -6740 53582 -6688
rect 53634 -6740 53644 -6688
rect 53767 -6740 53777 -6688
rect 53829 -6740 53839 -6688
rect 53957 -6740 53967 -6688
rect 54019 -6740 54029 -6688
rect 54148 -6740 54158 -6688
rect 54210 -6740 54220 -6688
rect 54340 -6740 54350 -6688
rect 54402 -6740 54412 -6688
rect 54533 -6739 54543 -6687
rect 54595 -6739 54605 -6687
rect 54725 -6740 54735 -6688
rect 54787 -6740 54797 -6688
rect 54917 -6740 54927 -6688
rect 54979 -6740 54989 -6688
rect 55110 -6740 55120 -6688
rect 55172 -6740 55182 -6688
rect 55301 -6739 55311 -6687
rect 55363 -6739 55373 -6687
rect 55493 -6740 55503 -6688
rect 55555 -6740 55565 -6688
rect 55685 -6739 55695 -6687
rect 55747 -6739 55757 -6687
rect 55877 -6739 55887 -6687
rect 55939 -6739 55949 -6687
rect 56068 -6740 56078 -6688
rect 56130 -6740 56140 -6688
rect 56261 -6739 56271 -6687
rect 56323 -6739 56333 -6687
rect 56453 -6739 56463 -6687
rect 56515 -6739 56525 -6687
rect 56647 -6740 56657 -6688
rect 56709 -6740 56719 -6688
rect 56838 -6741 56848 -6689
rect 56900 -6741 56910 -6689
rect 57027 -6740 57037 -6688
rect 57089 -6740 57099 -6688
rect 57220 -6740 57230 -6688
rect 57282 -6740 57292 -6688
rect 57413 -6740 57423 -6688
rect 57475 -6740 57485 -6688
rect 57604 -6739 57614 -6687
rect 57666 -6739 57676 -6687
rect 57795 -6739 57805 -6687
rect 57857 -6739 57867 -6687
rect 51940 -6880 51950 -6828
rect 52002 -6880 52012 -6828
rect 52132 -6880 52142 -6828
rect 52194 -6880 52204 -6828
rect 52325 -6880 52335 -6828
rect 52387 -6880 52397 -6828
rect 52517 -6880 52527 -6828
rect 52579 -6880 52589 -6828
rect 52710 -6880 52720 -6828
rect 52772 -6880 52782 -6828
rect 52902 -6879 52912 -6827
rect 52964 -6879 52974 -6827
rect 53093 -6880 53103 -6828
rect 53155 -6880 53165 -6828
rect 53285 -6880 53295 -6828
rect 53347 -6880 53357 -6828
rect 53477 -6879 53487 -6827
rect 53539 -6879 53549 -6827
rect 53669 -6879 53679 -6827
rect 53731 -6879 53741 -6827
rect 53861 -6880 53871 -6828
rect 53923 -6880 53933 -6828
rect 54053 -6879 54063 -6827
rect 54115 -6879 54125 -6827
rect 54245 -6880 54255 -6828
rect 54307 -6880 54317 -6828
rect 54436 -6879 54446 -6827
rect 54498 -6879 54508 -6827
rect 54630 -6880 54640 -6828
rect 54692 -6880 54702 -6828
rect 54820 -6880 54830 -6828
rect 54882 -6880 54892 -6828
rect 55012 -6880 55022 -6828
rect 55074 -6880 55084 -6828
rect 55205 -6880 55215 -6828
rect 55267 -6880 55277 -6828
rect 55396 -6880 55406 -6828
rect 55458 -6880 55468 -6828
rect 55589 -6879 55599 -6827
rect 55651 -6879 55661 -6827
rect 55782 -6880 55792 -6828
rect 55844 -6880 55854 -6828
rect 55973 -6880 55983 -6828
rect 56035 -6880 56045 -6828
rect 56166 -6880 56176 -6828
rect 56228 -6880 56238 -6828
rect 56356 -6880 56366 -6828
rect 56418 -6880 56428 -6828
rect 56550 -6879 56560 -6827
rect 56612 -6879 56622 -6827
rect 56739 -6880 56749 -6828
rect 56801 -6880 56811 -6828
rect 56932 -6880 56942 -6828
rect 56994 -6880 57004 -6828
rect 57125 -6880 57135 -6828
rect 57187 -6880 57197 -6828
rect 57315 -6880 57325 -6828
rect 57377 -6880 57387 -6828
rect 57508 -6879 57518 -6827
rect 57570 -6879 57580 -6827
rect 57697 -6879 57707 -6827
rect 57759 -6879 57769 -6827
rect 57900 -6920 57930 -6640
rect 51874 -6950 57930 -6920
rect 58070 -6640 64118 -6610
rect 58070 -6920 58100 -6640
rect 58226 -6740 58236 -6688
rect 58288 -6740 58298 -6688
rect 58416 -6739 58426 -6687
rect 58478 -6739 58488 -6687
rect 58608 -6738 58618 -6686
rect 58670 -6738 58680 -6686
rect 58799 -6738 58809 -6686
rect 58861 -6738 58871 -6686
rect 58993 -6738 59003 -6686
rect 59055 -6738 59065 -6686
rect 59183 -6739 59193 -6687
rect 59245 -6739 59255 -6687
rect 59377 -6738 59387 -6686
rect 59439 -6738 59449 -6686
rect 59569 -6738 59579 -6686
rect 59631 -6738 59641 -6686
rect 59760 -6739 59770 -6687
rect 59822 -6739 59832 -6687
rect 59955 -6739 59965 -6687
rect 60017 -6739 60027 -6687
rect 60145 -6739 60155 -6687
rect 60207 -6739 60217 -6687
rect 60336 -6739 60346 -6687
rect 60398 -6739 60408 -6687
rect 60528 -6739 60538 -6687
rect 60590 -6739 60600 -6687
rect 60721 -6738 60731 -6686
rect 60783 -6738 60793 -6686
rect 60913 -6739 60923 -6687
rect 60975 -6739 60985 -6687
rect 61105 -6739 61115 -6687
rect 61167 -6739 61177 -6687
rect 61298 -6739 61308 -6687
rect 61360 -6739 61370 -6687
rect 61489 -6738 61499 -6686
rect 61551 -6738 61561 -6686
rect 61681 -6739 61691 -6687
rect 61743 -6739 61753 -6687
rect 61873 -6738 61883 -6686
rect 61935 -6738 61945 -6686
rect 62065 -6738 62075 -6686
rect 62127 -6738 62137 -6686
rect 62256 -6739 62266 -6687
rect 62318 -6739 62328 -6687
rect 62449 -6738 62459 -6686
rect 62511 -6738 62521 -6686
rect 62641 -6738 62651 -6686
rect 62703 -6738 62713 -6686
rect 62835 -6739 62845 -6687
rect 62897 -6739 62907 -6687
rect 63026 -6740 63036 -6688
rect 63088 -6740 63098 -6688
rect 63215 -6739 63225 -6687
rect 63277 -6739 63287 -6687
rect 63408 -6739 63418 -6687
rect 63470 -6739 63480 -6687
rect 63601 -6739 63611 -6687
rect 63663 -6739 63673 -6687
rect 63792 -6738 63802 -6686
rect 63854 -6738 63864 -6686
rect 63983 -6738 63993 -6686
rect 64045 -6738 64055 -6686
rect 58130 -6879 58138 -6827
rect 58190 -6879 58200 -6827
rect 58320 -6879 58330 -6827
rect 58382 -6879 58392 -6827
rect 58513 -6879 58523 -6827
rect 58575 -6879 58585 -6827
rect 58705 -6879 58715 -6827
rect 58767 -6879 58777 -6827
rect 58898 -6879 58908 -6827
rect 58960 -6879 58970 -6827
rect 59090 -6878 59100 -6826
rect 59152 -6878 59162 -6826
rect 59281 -6879 59291 -6827
rect 59343 -6879 59353 -6827
rect 59473 -6879 59483 -6827
rect 59535 -6879 59545 -6827
rect 59665 -6878 59675 -6826
rect 59727 -6878 59737 -6826
rect 59857 -6878 59867 -6826
rect 59919 -6878 59929 -6826
rect 60049 -6879 60059 -6827
rect 60111 -6879 60121 -6827
rect 60241 -6878 60251 -6826
rect 60303 -6878 60313 -6826
rect 60433 -6879 60443 -6827
rect 60495 -6879 60505 -6827
rect 60624 -6878 60634 -6826
rect 60686 -6878 60696 -6826
rect 60818 -6879 60828 -6827
rect 60880 -6879 60890 -6827
rect 61008 -6879 61018 -6827
rect 61070 -6879 61080 -6827
rect 61200 -6879 61210 -6827
rect 61262 -6879 61272 -6827
rect 61393 -6879 61403 -6827
rect 61455 -6879 61465 -6827
rect 61584 -6879 61594 -6827
rect 61646 -6879 61656 -6827
rect 61777 -6878 61787 -6826
rect 61839 -6878 61849 -6826
rect 61970 -6879 61980 -6827
rect 62032 -6879 62042 -6827
rect 62161 -6879 62171 -6827
rect 62223 -6879 62233 -6827
rect 62354 -6879 62364 -6827
rect 62416 -6879 62426 -6827
rect 62544 -6879 62554 -6827
rect 62606 -6879 62616 -6827
rect 62738 -6878 62748 -6826
rect 62800 -6878 62810 -6826
rect 62927 -6879 62937 -6827
rect 62989 -6879 62999 -6827
rect 63120 -6879 63130 -6827
rect 63182 -6879 63192 -6827
rect 63313 -6879 63323 -6827
rect 63375 -6879 63385 -6827
rect 63503 -6879 63513 -6827
rect 63565 -6879 63575 -6827
rect 63696 -6878 63706 -6826
rect 63758 -6878 63768 -6826
rect 63885 -6878 63895 -6826
rect 63947 -6878 63957 -6826
rect 64084 -6920 64118 -6640
rect 66902 -6902 66912 -6850
rect 66964 -6902 66974 -6850
rect 58070 -6944 64118 -6920
rect 58070 -6950 64114 -6944
rect 49890 -7260 66624 -7230
rect 49890 -7312 49920 -7260
rect 49672 -7350 49920 -7312
rect 49672 -7584 49724 -7350
rect 49890 -7540 49920 -7350
rect 50077 -7354 50087 -7302
rect 50139 -7354 50149 -7302
rect 50267 -7353 50277 -7301
rect 50329 -7353 50339 -7301
rect 50460 -7356 50470 -7304
rect 50522 -7356 50532 -7304
rect 50652 -7351 50662 -7299
rect 50714 -7351 50724 -7299
rect 50844 -7355 50854 -7303
rect 50906 -7355 50916 -7303
rect 51036 -7350 51046 -7298
rect 51098 -7350 51108 -7298
rect 51228 -7351 51238 -7299
rect 51290 -7351 51300 -7299
rect 51418 -7350 51428 -7298
rect 51480 -7350 51490 -7298
rect 51612 -7361 51622 -7309
rect 51674 -7361 51684 -7309
rect 51801 -7359 51811 -7307
rect 51863 -7359 51873 -7307
rect 51991 -7359 52001 -7307
rect 52053 -7359 52063 -7307
rect 52190 -7360 52200 -7308
rect 52252 -7360 52262 -7308
rect 52382 -7359 52392 -7307
rect 52444 -7359 52454 -7307
rect 52572 -7360 52582 -7308
rect 52634 -7360 52644 -7308
rect 52764 -7353 52774 -7301
rect 52826 -7353 52836 -7301
rect 52956 -7303 53028 -7298
rect 52956 -7355 52966 -7303
rect 53018 -7355 53028 -7303
rect 53149 -7354 53159 -7302
rect 53211 -7354 53221 -7302
rect 53341 -7352 53351 -7300
rect 53403 -7352 53413 -7300
rect 53532 -7352 53542 -7300
rect 53594 -7352 53604 -7300
rect 53726 -7357 53736 -7305
rect 53788 -7357 53798 -7305
rect 53917 -7353 53927 -7301
rect 53979 -7353 53989 -7301
rect 54109 -7349 54119 -7297
rect 54171 -7349 54181 -7297
rect 54302 -7353 54312 -7301
rect 54364 -7353 54374 -7301
rect 54494 -7353 54504 -7301
rect 54556 -7353 54566 -7301
rect 54687 -7354 54697 -7302
rect 54749 -7354 54759 -7302
rect 54879 -7352 54889 -7300
rect 54941 -7352 54951 -7300
rect 55070 -7351 55080 -7299
rect 55132 -7351 55142 -7299
rect 55261 -7350 55271 -7298
rect 55323 -7350 55333 -7298
rect 55454 -7350 55464 -7298
rect 55516 -7350 55526 -7298
rect 55645 -7359 55655 -7307
rect 55707 -7359 55717 -7307
rect 55836 -7360 55846 -7308
rect 55898 -7360 55908 -7308
rect 56026 -7361 56036 -7309
rect 56088 -7361 56098 -7309
rect 56220 -7365 56230 -7313
rect 56282 -7365 56292 -7313
rect 56412 -7367 56422 -7315
rect 56474 -7367 56484 -7315
rect 56606 -7366 56616 -7314
rect 56668 -7366 56678 -7314
rect 56798 -7363 56808 -7311
rect 56860 -7363 56870 -7311
rect 56987 -7360 56997 -7308
rect 57049 -7360 57059 -7308
rect 57181 -7358 57191 -7306
rect 57243 -7358 57253 -7306
rect 57374 -7359 57384 -7307
rect 57436 -7359 57446 -7307
rect 57567 -7360 57577 -7308
rect 57629 -7360 57639 -7308
rect 57756 -7360 57766 -7308
rect 57818 -7360 57828 -7308
rect 57949 -7360 57959 -7308
rect 58011 -7360 58021 -7308
rect 58141 -7360 58151 -7308
rect 58203 -7360 58213 -7308
rect 58332 -7360 58342 -7308
rect 58394 -7360 58404 -7308
rect 58525 -7360 58535 -7308
rect 58587 -7360 58597 -7308
rect 58716 -7359 58726 -7307
rect 58778 -7359 58788 -7307
rect 58911 -7360 58921 -7308
rect 58973 -7360 58983 -7308
rect 59100 -7360 59110 -7308
rect 59162 -7360 59172 -7308
rect 59293 -7360 59303 -7308
rect 59355 -7360 59365 -7308
rect 59485 -7360 59495 -7308
rect 59547 -7360 59557 -7308
rect 59676 -7360 59686 -7308
rect 59738 -7360 59748 -7308
rect 59868 -7360 59878 -7308
rect 59930 -7360 59940 -7308
rect 60061 -7360 60071 -7308
rect 60123 -7360 60133 -7308
rect 60250 -7361 60260 -7309
rect 60312 -7361 60322 -7309
rect 60444 -7360 60454 -7308
rect 60506 -7360 60516 -7308
rect 60635 -7360 60645 -7308
rect 60697 -7360 60707 -7308
rect 60828 -7360 60838 -7308
rect 60890 -7360 60900 -7308
rect 61020 -7360 61030 -7308
rect 61082 -7360 61092 -7308
rect 61212 -7361 61222 -7309
rect 61274 -7361 61284 -7309
rect 61405 -7359 61415 -7307
rect 61467 -7359 61477 -7307
rect 61595 -7359 61605 -7307
rect 61657 -7359 61667 -7307
rect 61788 -7361 61798 -7309
rect 61850 -7361 61860 -7309
rect 61980 -7360 61990 -7308
rect 62042 -7360 62052 -7308
rect 62173 -7359 62183 -7307
rect 62235 -7359 62245 -7307
rect 62364 -7359 62374 -7307
rect 62426 -7359 62436 -7307
rect 62556 -7360 62566 -7308
rect 62618 -7360 62628 -7308
rect 62747 -7360 62757 -7308
rect 62809 -7360 62819 -7308
rect 62939 -7360 62949 -7308
rect 63001 -7360 63011 -7308
rect 63133 -7359 63143 -7307
rect 63195 -7359 63205 -7307
rect 63325 -7360 63335 -7308
rect 63387 -7360 63397 -7308
rect 63515 -7361 63525 -7309
rect 63577 -7361 63587 -7309
rect 63706 -7362 63716 -7310
rect 63768 -7362 63778 -7310
rect 63899 -7360 63909 -7308
rect 63961 -7360 63971 -7308
rect 64092 -7359 64102 -7307
rect 64154 -7359 64164 -7307
rect 64285 -7360 64295 -7308
rect 64347 -7360 64357 -7308
rect 64476 -7360 64486 -7308
rect 64538 -7360 64548 -7308
rect 64667 -7360 64677 -7308
rect 64729 -7360 64739 -7308
rect 64860 -7360 64870 -7308
rect 64922 -7360 64932 -7308
rect 65053 -7360 65063 -7308
rect 65115 -7360 65125 -7308
rect 65244 -7360 65254 -7308
rect 65306 -7360 65316 -7308
rect 65435 -7359 65445 -7307
rect 65497 -7359 65507 -7307
rect 65626 -7359 65636 -7307
rect 65688 -7359 65698 -7307
rect 65819 -7360 65829 -7308
rect 65881 -7360 65891 -7308
rect 66013 -7360 66023 -7308
rect 66075 -7360 66085 -7308
rect 66201 -7361 66211 -7309
rect 66263 -7361 66273 -7309
rect 66395 -7369 66405 -7317
rect 66457 -7369 66467 -7317
rect 49981 -7497 49991 -7445
rect 50043 -7497 50053 -7445
rect 50172 -7499 50182 -7447
rect 50234 -7499 50244 -7447
rect 50364 -7498 50374 -7446
rect 50426 -7498 50436 -7446
rect 50556 -7501 50566 -7449
rect 50618 -7501 50628 -7449
rect 50750 -7500 50760 -7448
rect 50812 -7500 50822 -7448
rect 50940 -7500 50950 -7448
rect 51002 -7500 51012 -7448
rect 51135 -7498 51145 -7446
rect 51197 -7498 51207 -7446
rect 51326 -7497 51336 -7445
rect 51388 -7497 51398 -7445
rect 51521 -7499 51531 -7447
rect 51583 -7499 51593 -7447
rect 51711 -7499 51721 -7447
rect 51773 -7499 51783 -7447
rect 51901 -7498 51911 -7446
rect 51963 -7498 51973 -7446
rect 52094 -7497 52104 -7445
rect 52156 -7497 52166 -7445
rect 52285 -7497 52295 -7445
rect 52347 -7497 52357 -7445
rect 52481 -7499 52491 -7447
rect 52543 -7499 52553 -7447
rect 52670 -7499 52680 -7447
rect 52732 -7499 52742 -7447
rect 52864 -7499 52874 -7447
rect 52926 -7499 52936 -7447
rect 53053 -7499 53063 -7447
rect 53115 -7499 53125 -7447
rect 53245 -7500 53255 -7448
rect 53307 -7500 53317 -7448
rect 53438 -7500 53448 -7448
rect 53500 -7500 53510 -7448
rect 53629 -7500 53639 -7448
rect 53691 -7500 53701 -7448
rect 53821 -7499 53831 -7447
rect 53883 -7499 53893 -7447
rect 54013 -7500 54023 -7448
rect 54075 -7500 54085 -7448
rect 54206 -7500 54216 -7448
rect 54268 -7500 54278 -7448
rect 54397 -7500 54407 -7448
rect 54459 -7500 54469 -7448
rect 54589 -7499 54599 -7447
rect 54651 -7499 54661 -7447
rect 54782 -7500 54792 -7448
rect 54844 -7500 54854 -7448
rect 54974 -7500 54984 -7448
rect 55036 -7500 55046 -7448
rect 55165 -7500 55175 -7448
rect 55227 -7500 55237 -7448
rect 55356 -7500 55366 -7448
rect 55418 -7500 55428 -7448
rect 55548 -7500 55558 -7448
rect 55610 -7500 55620 -7448
rect 55741 -7499 55751 -7447
rect 55803 -7499 55813 -7447
rect 55932 -7499 55942 -7447
rect 55994 -7499 56004 -7447
rect 56126 -7500 56136 -7448
rect 56188 -7500 56198 -7448
rect 56318 -7500 56328 -7448
rect 56380 -7500 56390 -7448
rect 56510 -7500 56520 -7448
rect 56572 -7500 56582 -7448
rect 56702 -7500 56712 -7448
rect 56764 -7500 56774 -7448
rect 56894 -7500 56904 -7448
rect 56956 -7500 56966 -7448
rect 57086 -7500 57096 -7448
rect 57148 -7500 57158 -7448
rect 57278 -7500 57288 -7448
rect 57340 -7500 57350 -7448
rect 57469 -7500 57479 -7448
rect 57531 -7500 57541 -7448
rect 57661 -7500 57671 -7448
rect 57723 -7500 57733 -7448
rect 57854 -7500 57864 -7448
rect 57916 -7500 57926 -7448
rect 58046 -7500 58056 -7448
rect 58108 -7500 58118 -7448
rect 58238 -7500 58248 -7448
rect 58300 -7500 58310 -7448
rect 58429 -7500 58439 -7448
rect 58491 -7500 58501 -7448
rect 58621 -7500 58631 -7448
rect 58683 -7500 58693 -7448
rect 58812 -7500 58822 -7448
rect 58874 -7500 58884 -7448
rect 59003 -7500 59013 -7448
rect 59065 -7500 59075 -7448
rect 59197 -7500 59207 -7448
rect 59259 -7500 59269 -7448
rect 59389 -7500 59399 -7448
rect 59451 -7500 59461 -7448
rect 59582 -7499 59592 -7447
rect 59644 -7499 59654 -7447
rect 59773 -7500 59783 -7448
rect 59835 -7500 59845 -7448
rect 59965 -7500 59975 -7448
rect 60027 -7500 60037 -7448
rect 60158 -7500 60168 -7448
rect 60220 -7500 60230 -7448
rect 60350 -7500 60360 -7448
rect 60412 -7500 60422 -7448
rect 60543 -7499 60553 -7447
rect 60605 -7499 60615 -7447
rect 60734 -7500 60744 -7448
rect 60796 -7500 60806 -7448
rect 60926 -7500 60936 -7448
rect 60988 -7500 60998 -7448
rect 61117 -7500 61127 -7448
rect 61179 -7500 61189 -7448
rect 61309 -7500 61319 -7448
rect 61371 -7500 61381 -7448
rect 61501 -7500 61511 -7448
rect 61563 -7500 61573 -7448
rect 61694 -7500 61704 -7448
rect 61756 -7500 61766 -7448
rect 61885 -7500 61895 -7448
rect 61947 -7500 61957 -7448
rect 62077 -7500 62087 -7448
rect 62139 -7500 62149 -7448
rect 62269 -7499 62279 -7447
rect 62331 -7499 62341 -7447
rect 62461 -7500 62471 -7448
rect 62523 -7500 62533 -7448
rect 62651 -7500 62661 -7448
rect 62713 -7500 62723 -7448
rect 62845 -7500 62855 -7448
rect 62907 -7500 62917 -7448
rect 63037 -7499 63047 -7447
rect 63099 -7499 63109 -7447
rect 63228 -7500 63238 -7448
rect 63290 -7500 63300 -7448
rect 63421 -7500 63431 -7448
rect 63483 -7500 63493 -7448
rect 63612 -7499 63622 -7447
rect 63674 -7499 63684 -7447
rect 63804 -7500 63814 -7448
rect 63866 -7500 63876 -7448
rect 63995 -7500 64005 -7448
rect 64057 -7500 64067 -7448
rect 64189 -7499 64199 -7447
rect 64251 -7499 64261 -7447
rect 64380 -7500 64390 -7448
rect 64442 -7500 64452 -7448
rect 64572 -7500 64582 -7448
rect 64634 -7500 64644 -7448
rect 64764 -7500 64774 -7448
rect 64826 -7500 64836 -7448
rect 64956 -7500 64966 -7448
rect 65018 -7500 65028 -7448
rect 65149 -7500 65159 -7448
rect 65211 -7500 65221 -7448
rect 65340 -7500 65350 -7448
rect 65402 -7500 65412 -7448
rect 65533 -7499 65543 -7447
rect 65595 -7499 65605 -7447
rect 65724 -7500 65734 -7448
rect 65786 -7500 65796 -7448
rect 65917 -7500 65927 -7448
rect 65979 -7500 65989 -7448
rect 66108 -7500 66118 -7448
rect 66170 -7500 66180 -7448
rect 66299 -7498 66309 -7446
rect 66361 -7498 66371 -7446
rect 66494 -7500 66504 -7448
rect 66556 -7500 66566 -7448
rect 66594 -7540 66624 -7260
rect 66912 -7270 66974 -6902
rect 68006 -7234 68368 -6644
rect 68006 -7270 68374 -7234
rect 66912 -7334 68374 -7270
rect 66932 -7338 68374 -7334
rect 49890 -7570 66624 -7540
rect 68006 -7640 68374 -7338
rect 68368 -7642 68374 -7640
rect 49928 -7664 66600 -7658
rect 49928 -7692 49940 -7664
rect 48262 -7706 48458 -7700
rect 48262 -7764 48274 -7706
rect 48446 -7764 48458 -7706
rect 49524 -7752 49940 -7692
rect 49928 -7756 49940 -7752
rect 66588 -7756 66600 -7664
rect 49928 -7762 66600 -7756
rect 68108 -7710 68304 -7704
rect 48262 -7770 48458 -7764
rect 68108 -7768 68120 -7710
rect 68292 -7768 68304 -7710
rect 68914 -7756 68924 -6672
rect 69290 -7756 69300 -6672
rect 68108 -7774 68304 -7768
<< via1 >>
rect 47254 -7752 47614 -6678
rect 49436 -6924 49488 -6872
rect 52048 -6741 52100 -6689
rect 52238 -6740 52290 -6688
rect 52430 -6739 52482 -6687
rect 52621 -6739 52673 -6687
rect 52815 -6739 52867 -6687
rect 53005 -6740 53057 -6688
rect 53199 -6739 53251 -6687
rect 53391 -6739 53443 -6687
rect 53582 -6740 53634 -6688
rect 53777 -6740 53829 -6688
rect 53967 -6740 54019 -6688
rect 54158 -6740 54210 -6688
rect 54350 -6740 54402 -6688
rect 54543 -6739 54595 -6687
rect 54735 -6740 54787 -6688
rect 54927 -6740 54979 -6688
rect 55120 -6740 55172 -6688
rect 55311 -6739 55363 -6687
rect 55503 -6740 55555 -6688
rect 55695 -6739 55747 -6687
rect 55887 -6739 55939 -6687
rect 56078 -6740 56130 -6688
rect 56271 -6739 56323 -6687
rect 56463 -6739 56515 -6687
rect 56657 -6740 56709 -6688
rect 56848 -6741 56900 -6689
rect 57037 -6740 57089 -6688
rect 57230 -6740 57282 -6688
rect 57423 -6740 57475 -6688
rect 57614 -6739 57666 -6687
rect 57805 -6739 57857 -6687
rect 51950 -6880 52002 -6828
rect 52142 -6880 52194 -6828
rect 52335 -6880 52387 -6828
rect 52527 -6880 52579 -6828
rect 52720 -6880 52772 -6828
rect 52912 -6879 52964 -6827
rect 53103 -6880 53155 -6828
rect 53295 -6880 53347 -6828
rect 53487 -6879 53539 -6827
rect 53679 -6879 53731 -6827
rect 53871 -6880 53923 -6828
rect 54063 -6879 54115 -6827
rect 54255 -6880 54307 -6828
rect 54446 -6879 54498 -6827
rect 54640 -6880 54692 -6828
rect 54830 -6880 54882 -6828
rect 55022 -6880 55074 -6828
rect 55215 -6880 55267 -6828
rect 55406 -6880 55458 -6828
rect 55599 -6879 55651 -6827
rect 55792 -6880 55844 -6828
rect 55983 -6880 56035 -6828
rect 56176 -6880 56228 -6828
rect 56366 -6880 56418 -6828
rect 56560 -6879 56612 -6827
rect 56749 -6880 56801 -6828
rect 56942 -6880 56994 -6828
rect 57135 -6880 57187 -6828
rect 57325 -6880 57377 -6828
rect 57518 -6879 57570 -6827
rect 57707 -6879 57759 -6827
rect 58236 -6740 58288 -6688
rect 58426 -6739 58478 -6687
rect 58618 -6738 58670 -6686
rect 58809 -6738 58861 -6686
rect 59003 -6738 59055 -6686
rect 59193 -6739 59245 -6687
rect 59387 -6738 59439 -6686
rect 59579 -6738 59631 -6686
rect 59770 -6739 59822 -6687
rect 59965 -6739 60017 -6687
rect 60155 -6739 60207 -6687
rect 60346 -6739 60398 -6687
rect 60538 -6739 60590 -6687
rect 60731 -6738 60783 -6686
rect 60923 -6739 60975 -6687
rect 61115 -6739 61167 -6687
rect 61308 -6739 61360 -6687
rect 61499 -6738 61551 -6686
rect 61691 -6739 61743 -6687
rect 61883 -6738 61935 -6686
rect 62075 -6738 62127 -6686
rect 62266 -6739 62318 -6687
rect 62459 -6738 62511 -6686
rect 62651 -6738 62703 -6686
rect 62845 -6739 62897 -6687
rect 63036 -6740 63088 -6688
rect 63225 -6739 63277 -6687
rect 63418 -6739 63470 -6687
rect 63611 -6739 63663 -6687
rect 63802 -6738 63854 -6686
rect 63993 -6738 64045 -6686
rect 58138 -6879 58190 -6827
rect 58330 -6879 58382 -6827
rect 58523 -6879 58575 -6827
rect 58715 -6879 58767 -6827
rect 58908 -6879 58960 -6827
rect 59100 -6878 59152 -6826
rect 59291 -6879 59343 -6827
rect 59483 -6879 59535 -6827
rect 59675 -6878 59727 -6826
rect 59867 -6878 59919 -6826
rect 60059 -6879 60111 -6827
rect 60251 -6878 60303 -6826
rect 60443 -6879 60495 -6827
rect 60634 -6878 60686 -6826
rect 60828 -6879 60880 -6827
rect 61018 -6879 61070 -6827
rect 61210 -6879 61262 -6827
rect 61403 -6879 61455 -6827
rect 61594 -6879 61646 -6827
rect 61787 -6878 61839 -6826
rect 61980 -6879 62032 -6827
rect 62171 -6879 62223 -6827
rect 62364 -6879 62416 -6827
rect 62554 -6879 62606 -6827
rect 62748 -6878 62800 -6826
rect 62937 -6879 62989 -6827
rect 63130 -6879 63182 -6827
rect 63323 -6879 63375 -6827
rect 63513 -6879 63565 -6827
rect 63706 -6878 63758 -6826
rect 63895 -6878 63947 -6826
rect 66912 -6902 66964 -6850
rect 50087 -7354 50139 -7302
rect 50277 -7353 50329 -7301
rect 50470 -7356 50522 -7304
rect 50662 -7351 50714 -7299
rect 50854 -7355 50906 -7303
rect 51046 -7350 51098 -7298
rect 51238 -7351 51290 -7299
rect 51428 -7350 51480 -7298
rect 51622 -7361 51674 -7309
rect 51811 -7359 51863 -7307
rect 52001 -7359 52053 -7307
rect 52200 -7360 52252 -7308
rect 52392 -7359 52444 -7307
rect 52582 -7360 52634 -7308
rect 52774 -7353 52826 -7301
rect 52966 -7355 53018 -7303
rect 53159 -7354 53211 -7302
rect 53351 -7352 53403 -7300
rect 53542 -7352 53594 -7300
rect 53736 -7357 53788 -7305
rect 53927 -7353 53979 -7301
rect 54119 -7349 54171 -7297
rect 54312 -7353 54364 -7301
rect 54504 -7353 54556 -7301
rect 54697 -7354 54749 -7302
rect 54889 -7352 54941 -7300
rect 55080 -7351 55132 -7299
rect 55271 -7350 55323 -7298
rect 55464 -7350 55516 -7298
rect 55655 -7359 55707 -7307
rect 55846 -7360 55898 -7308
rect 56036 -7361 56088 -7309
rect 56230 -7365 56282 -7313
rect 56422 -7367 56474 -7315
rect 56616 -7366 56668 -7314
rect 56808 -7363 56860 -7311
rect 56997 -7360 57049 -7308
rect 57191 -7358 57243 -7306
rect 57384 -7359 57436 -7307
rect 57577 -7360 57629 -7308
rect 57766 -7360 57818 -7308
rect 57959 -7360 58011 -7308
rect 58151 -7360 58203 -7308
rect 58342 -7360 58394 -7308
rect 58535 -7360 58587 -7308
rect 58726 -7359 58778 -7307
rect 58921 -7360 58973 -7308
rect 59110 -7360 59162 -7308
rect 59303 -7360 59355 -7308
rect 59495 -7360 59547 -7308
rect 59686 -7360 59738 -7308
rect 59878 -7360 59930 -7308
rect 60071 -7360 60123 -7308
rect 60260 -7361 60312 -7309
rect 60454 -7360 60506 -7308
rect 60645 -7360 60697 -7308
rect 60838 -7360 60890 -7308
rect 61030 -7360 61082 -7308
rect 61222 -7361 61274 -7309
rect 61415 -7359 61467 -7307
rect 61605 -7359 61657 -7307
rect 61798 -7361 61850 -7309
rect 61990 -7360 62042 -7308
rect 62183 -7359 62235 -7307
rect 62374 -7359 62426 -7307
rect 62566 -7360 62618 -7308
rect 62757 -7360 62809 -7308
rect 62949 -7360 63001 -7308
rect 63143 -7359 63195 -7307
rect 63335 -7360 63387 -7308
rect 63525 -7361 63577 -7309
rect 63716 -7362 63768 -7310
rect 63909 -7360 63961 -7308
rect 64102 -7359 64154 -7307
rect 64295 -7360 64347 -7308
rect 64486 -7360 64538 -7308
rect 64677 -7360 64729 -7308
rect 64870 -7360 64922 -7308
rect 65063 -7360 65115 -7308
rect 65254 -7360 65306 -7308
rect 65445 -7359 65497 -7307
rect 65636 -7359 65688 -7307
rect 65829 -7360 65881 -7308
rect 66023 -7360 66075 -7308
rect 66211 -7361 66263 -7309
rect 66405 -7369 66457 -7317
rect 49991 -7497 50043 -7445
rect 50182 -7499 50234 -7447
rect 50374 -7498 50426 -7446
rect 50566 -7501 50618 -7449
rect 50760 -7500 50812 -7448
rect 50950 -7500 51002 -7448
rect 51145 -7498 51197 -7446
rect 51336 -7497 51388 -7445
rect 51531 -7499 51583 -7447
rect 51721 -7499 51773 -7447
rect 51911 -7498 51963 -7446
rect 52104 -7497 52156 -7445
rect 52295 -7497 52347 -7445
rect 52491 -7499 52543 -7447
rect 52680 -7499 52732 -7447
rect 52874 -7499 52926 -7447
rect 53063 -7499 53115 -7447
rect 53255 -7500 53307 -7448
rect 53448 -7500 53500 -7448
rect 53639 -7500 53691 -7448
rect 53831 -7499 53883 -7447
rect 54023 -7500 54075 -7448
rect 54216 -7500 54268 -7448
rect 54407 -7500 54459 -7448
rect 54599 -7499 54651 -7447
rect 54792 -7500 54844 -7448
rect 54984 -7500 55036 -7448
rect 55175 -7500 55227 -7448
rect 55366 -7500 55418 -7448
rect 55558 -7500 55610 -7448
rect 55751 -7499 55803 -7447
rect 55942 -7499 55994 -7447
rect 56136 -7500 56188 -7448
rect 56328 -7500 56380 -7448
rect 56520 -7500 56572 -7448
rect 56712 -7500 56764 -7448
rect 56904 -7500 56956 -7448
rect 57096 -7500 57148 -7448
rect 57288 -7500 57340 -7448
rect 57479 -7500 57531 -7448
rect 57671 -7500 57723 -7448
rect 57864 -7500 57916 -7448
rect 58056 -7500 58108 -7448
rect 58248 -7500 58300 -7448
rect 58439 -7500 58491 -7448
rect 58631 -7500 58683 -7448
rect 58822 -7500 58874 -7448
rect 59013 -7500 59065 -7448
rect 59207 -7500 59259 -7448
rect 59399 -7500 59451 -7448
rect 59592 -7499 59644 -7447
rect 59783 -7500 59835 -7448
rect 59975 -7500 60027 -7448
rect 60168 -7500 60220 -7448
rect 60360 -7500 60412 -7448
rect 60553 -7499 60605 -7447
rect 60744 -7500 60796 -7448
rect 60936 -7500 60988 -7448
rect 61127 -7500 61179 -7448
rect 61319 -7500 61371 -7448
rect 61511 -7500 61563 -7448
rect 61704 -7500 61756 -7448
rect 61895 -7500 61947 -7448
rect 62087 -7500 62139 -7448
rect 62279 -7499 62331 -7447
rect 62471 -7500 62523 -7448
rect 62661 -7500 62713 -7448
rect 62855 -7500 62907 -7448
rect 63047 -7499 63099 -7447
rect 63238 -7500 63290 -7448
rect 63431 -7500 63483 -7448
rect 63622 -7499 63674 -7447
rect 63814 -7500 63866 -7448
rect 64005 -7500 64057 -7448
rect 64199 -7499 64251 -7447
rect 64390 -7500 64442 -7448
rect 64582 -7500 64634 -7448
rect 64774 -7500 64826 -7448
rect 64966 -7500 65018 -7448
rect 65159 -7500 65211 -7448
rect 65350 -7500 65402 -7448
rect 65543 -7499 65595 -7447
rect 65734 -7500 65786 -7448
rect 65927 -7500 65979 -7448
rect 66118 -7500 66170 -7448
rect 66309 -7498 66361 -7446
rect 66504 -7500 66556 -7448
rect 48274 -7764 48446 -7706
rect 49940 -7756 66588 -7664
rect 68120 -7768 68292 -7710
rect 68924 -7756 69290 -6672
<< metal2 >>
rect 47224 -6678 47652 -6366
rect 47224 -7752 47254 -6678
rect 47614 -7752 47652 -6678
rect 52040 -6680 52100 -6434
rect 52238 -6680 52290 -6678
rect 52430 -6680 52482 -6677
rect 52621 -6680 52673 -6677
rect 52815 -6680 52867 -6677
rect 53005 -6680 53057 -6678
rect 53199 -6680 53251 -6677
rect 53391 -6680 53443 -6677
rect 53582 -6680 53634 -6678
rect 53777 -6680 53829 -6678
rect 53967 -6680 54019 -6678
rect 54158 -6680 54210 -6678
rect 54350 -6680 54402 -6678
rect 54543 -6680 54595 -6677
rect 54735 -6680 54787 -6678
rect 54927 -6680 54979 -6678
rect 55120 -6680 55172 -6678
rect 55311 -6680 55363 -6677
rect 55503 -6680 55555 -6678
rect 55695 -6680 55747 -6677
rect 55887 -6680 55939 -6677
rect 56078 -6680 56130 -6678
rect 56271 -6680 56323 -6677
rect 56463 -6680 56515 -6677
rect 56657 -6680 56709 -6678
rect 56848 -6680 56900 -6679
rect 57037 -6680 57089 -6678
rect 57230 -6680 57282 -6678
rect 57423 -6680 57475 -6678
rect 57614 -6680 57666 -6677
rect 57800 -6680 57860 -6388
rect 49440 -6687 57860 -6680
rect 49440 -6688 52430 -6687
rect 49440 -6689 52238 -6688
rect 49440 -6720 52048 -6689
rect 49440 -6862 49470 -6720
rect 52100 -6710 52238 -6689
rect 52048 -6751 52100 -6741
rect 52290 -6710 52430 -6688
rect 52238 -6750 52290 -6740
rect 52482 -6710 52621 -6687
rect 52430 -6749 52482 -6739
rect 52673 -6710 52815 -6687
rect 52621 -6749 52673 -6739
rect 52867 -6688 53199 -6687
rect 52867 -6710 53005 -6688
rect 52815 -6749 52867 -6739
rect 53057 -6710 53199 -6688
rect 53005 -6750 53057 -6740
rect 53251 -6710 53391 -6687
rect 53199 -6749 53251 -6739
rect 53443 -6688 54543 -6687
rect 53443 -6710 53582 -6688
rect 53391 -6749 53443 -6739
rect 53634 -6710 53777 -6688
rect 53582 -6750 53634 -6740
rect 53829 -6710 53967 -6688
rect 53777 -6750 53829 -6740
rect 54019 -6710 54158 -6688
rect 53967 -6750 54019 -6740
rect 54210 -6710 54350 -6688
rect 54158 -6750 54210 -6740
rect 54402 -6710 54543 -6688
rect 54350 -6750 54402 -6740
rect 54595 -6688 55311 -6687
rect 54595 -6710 54735 -6688
rect 54543 -6749 54595 -6739
rect 54787 -6710 54927 -6688
rect 54735 -6750 54787 -6740
rect 54979 -6710 55120 -6688
rect 54927 -6750 54979 -6740
rect 55172 -6710 55311 -6688
rect 55120 -6750 55172 -6740
rect 55363 -6688 55695 -6687
rect 55363 -6710 55503 -6688
rect 55311 -6749 55363 -6739
rect 55555 -6710 55695 -6688
rect 55503 -6750 55555 -6740
rect 55747 -6710 55887 -6687
rect 55695 -6749 55747 -6739
rect 55939 -6688 56271 -6687
rect 55939 -6710 56078 -6688
rect 55887 -6749 55939 -6739
rect 56130 -6710 56271 -6688
rect 56078 -6750 56130 -6740
rect 56323 -6710 56463 -6687
rect 56271 -6749 56323 -6739
rect 56515 -6688 57614 -6687
rect 56515 -6710 56657 -6688
rect 56463 -6749 56515 -6739
rect 56709 -6689 57037 -6688
rect 56709 -6710 56848 -6689
rect 56657 -6750 56709 -6740
rect 56900 -6710 57037 -6689
rect 56848 -6751 56900 -6741
rect 57089 -6710 57230 -6688
rect 57037 -6750 57089 -6740
rect 57282 -6710 57423 -6688
rect 57230 -6750 57282 -6740
rect 57475 -6710 57614 -6688
rect 57423 -6750 57475 -6740
rect 57666 -6710 57805 -6687
rect 57614 -6749 57666 -6739
rect 57857 -6690 57860 -6687
rect 58230 -6679 58290 -6398
rect 58426 -6679 58478 -6677
rect 58618 -6679 58670 -6676
rect 58809 -6679 58861 -6676
rect 59003 -6679 59055 -6676
rect 59193 -6679 59245 -6677
rect 59387 -6679 59439 -6676
rect 59579 -6679 59631 -6676
rect 59770 -6679 59822 -6677
rect 59965 -6679 60017 -6677
rect 60155 -6679 60207 -6677
rect 60346 -6679 60398 -6677
rect 60538 -6679 60590 -6677
rect 60731 -6679 60783 -6676
rect 60923 -6679 60975 -6677
rect 61115 -6679 61167 -6677
rect 61308 -6679 61360 -6677
rect 61499 -6679 61551 -6676
rect 61691 -6679 61743 -6677
rect 61883 -6679 61935 -6676
rect 62075 -6679 62127 -6676
rect 62266 -6679 62318 -6677
rect 62459 -6679 62511 -6676
rect 62651 -6679 62703 -6676
rect 62845 -6679 62897 -6677
rect 63036 -6679 63088 -6678
rect 63225 -6679 63277 -6677
rect 63418 -6679 63470 -6677
rect 63611 -6679 63663 -6677
rect 63802 -6679 63854 -6676
rect 63990 -6679 64050 -6366
rect 58230 -6680 64050 -6679
rect 68894 -6672 69326 -6366
rect 58230 -6686 66950 -6680
rect 58230 -6687 58618 -6686
rect 58230 -6688 58426 -6687
rect 58230 -6690 58236 -6688
rect 57805 -6749 57857 -6739
rect 58288 -6709 58426 -6688
rect 58236 -6750 58288 -6740
rect 58478 -6709 58618 -6687
rect 58426 -6749 58478 -6739
rect 58670 -6709 58809 -6686
rect 58618 -6748 58670 -6738
rect 58861 -6709 59003 -6686
rect 58809 -6748 58861 -6738
rect 59055 -6687 59387 -6686
rect 59055 -6709 59193 -6687
rect 59003 -6748 59055 -6738
rect 59245 -6709 59387 -6687
rect 59193 -6749 59245 -6739
rect 59439 -6709 59579 -6686
rect 59387 -6748 59439 -6738
rect 59631 -6687 60731 -6686
rect 59631 -6709 59770 -6687
rect 59579 -6748 59631 -6738
rect 59822 -6709 59965 -6687
rect 59770 -6749 59822 -6739
rect 60017 -6709 60155 -6687
rect 59965 -6749 60017 -6739
rect 60207 -6709 60346 -6687
rect 60155 -6749 60207 -6739
rect 60398 -6709 60538 -6687
rect 60346 -6749 60398 -6739
rect 60590 -6709 60731 -6687
rect 60538 -6749 60590 -6739
rect 60783 -6687 61499 -6686
rect 60783 -6709 60923 -6687
rect 60731 -6748 60783 -6738
rect 60975 -6709 61115 -6687
rect 60923 -6749 60975 -6739
rect 61167 -6709 61308 -6687
rect 61115 -6749 61167 -6739
rect 61360 -6709 61499 -6687
rect 61308 -6749 61360 -6739
rect 61551 -6687 61883 -6686
rect 61551 -6709 61691 -6687
rect 61499 -6748 61551 -6738
rect 61743 -6709 61883 -6687
rect 61691 -6749 61743 -6739
rect 61935 -6709 62075 -6686
rect 61883 -6748 61935 -6738
rect 62127 -6687 62459 -6686
rect 62127 -6709 62266 -6687
rect 62075 -6748 62127 -6738
rect 62318 -6709 62459 -6687
rect 62266 -6749 62318 -6739
rect 62511 -6709 62651 -6686
rect 62459 -6748 62511 -6738
rect 62703 -6687 63802 -6686
rect 62703 -6709 62845 -6687
rect 62651 -6748 62703 -6738
rect 62897 -6688 63225 -6687
rect 62897 -6709 63036 -6688
rect 62845 -6749 62897 -6739
rect 63088 -6709 63225 -6688
rect 63036 -6750 63088 -6740
rect 63277 -6709 63418 -6687
rect 63225 -6749 63277 -6739
rect 63470 -6709 63611 -6687
rect 63418 -6749 63470 -6739
rect 63663 -6709 63802 -6687
rect 63611 -6749 63663 -6739
rect 63854 -6709 63993 -6686
rect 63802 -6748 63854 -6738
rect 64045 -6710 66950 -6686
rect 63993 -6748 64045 -6738
rect 51950 -6826 63950 -6810
rect 51950 -6827 59100 -6826
rect 51950 -6828 52912 -6827
rect 49436 -6872 49488 -6862
rect 52002 -6880 52142 -6828
rect 52194 -6880 52335 -6828
rect 52387 -6880 52527 -6828
rect 52579 -6880 52720 -6828
rect 52772 -6879 52912 -6828
rect 52964 -6828 53487 -6827
rect 52964 -6879 53103 -6828
rect 52772 -6880 53103 -6879
rect 53155 -6880 53295 -6828
rect 53347 -6879 53487 -6828
rect 53539 -6879 53679 -6827
rect 53731 -6828 54063 -6827
rect 53731 -6879 53871 -6828
rect 53347 -6880 53871 -6879
rect 53923 -6879 54063 -6828
rect 54115 -6828 54446 -6827
rect 54115 -6879 54255 -6828
rect 53923 -6880 54255 -6879
rect 54307 -6879 54446 -6828
rect 54498 -6828 55599 -6827
rect 54498 -6879 54640 -6828
rect 54307 -6880 54640 -6879
rect 54692 -6880 54830 -6828
rect 54882 -6880 55022 -6828
rect 55074 -6880 55215 -6828
rect 55267 -6880 55406 -6828
rect 55458 -6879 55599 -6828
rect 55651 -6828 56560 -6827
rect 55651 -6879 55792 -6828
rect 55458 -6880 55792 -6879
rect 55844 -6880 55983 -6828
rect 56035 -6880 56176 -6828
rect 56228 -6880 56366 -6828
rect 56418 -6879 56560 -6828
rect 56612 -6828 57518 -6827
rect 56612 -6879 56749 -6828
rect 56418 -6880 56749 -6879
rect 56801 -6880 56942 -6828
rect 56994 -6880 57135 -6828
rect 57187 -6880 57325 -6828
rect 57377 -6879 57518 -6828
rect 57570 -6879 57707 -6827
rect 57759 -6879 58138 -6827
rect 58190 -6879 58330 -6827
rect 58382 -6879 58523 -6827
rect 58575 -6879 58715 -6827
rect 58767 -6879 58908 -6827
rect 58960 -6878 59100 -6827
rect 59152 -6827 59675 -6826
rect 59152 -6878 59291 -6827
rect 58960 -6879 59291 -6878
rect 59343 -6879 59483 -6827
rect 59535 -6878 59675 -6827
rect 59727 -6878 59867 -6826
rect 59919 -6827 60251 -6826
rect 59919 -6878 60059 -6827
rect 59535 -6879 60059 -6878
rect 60111 -6878 60251 -6827
rect 60303 -6827 60634 -6826
rect 60303 -6878 60443 -6827
rect 60111 -6879 60443 -6878
rect 60495 -6878 60634 -6827
rect 60686 -6827 61787 -6826
rect 60686 -6878 60828 -6827
rect 60495 -6879 60828 -6878
rect 60880 -6879 61018 -6827
rect 61070 -6879 61210 -6827
rect 61262 -6879 61403 -6827
rect 61455 -6879 61594 -6827
rect 61646 -6878 61787 -6827
rect 61839 -6827 62748 -6826
rect 61839 -6878 61980 -6827
rect 61646 -6879 61980 -6878
rect 62032 -6879 62171 -6827
rect 62223 -6879 62364 -6827
rect 62416 -6879 62554 -6827
rect 62606 -6878 62748 -6827
rect 62800 -6827 63706 -6826
rect 62800 -6878 62937 -6827
rect 62606 -6879 62937 -6878
rect 62989 -6879 63130 -6827
rect 63182 -6879 63323 -6827
rect 63375 -6879 63513 -6827
rect 63565 -6878 63706 -6827
rect 63758 -6878 63895 -6826
rect 63947 -6878 63950 -6826
rect 66920 -6840 66950 -6710
rect 63565 -6879 63950 -6878
rect 57377 -6880 63950 -6879
rect 51950 -6890 63950 -6880
rect 66912 -6850 66964 -6840
rect 49436 -6934 49488 -6924
rect 50087 -7300 50139 -7292
rect 50277 -7300 50329 -7291
rect 50470 -7300 50522 -7294
rect 50662 -7299 50714 -7289
rect 50087 -7301 50662 -7300
rect 50087 -7302 50277 -7301
rect 50139 -7330 50277 -7302
rect 50087 -7364 50139 -7354
rect 50329 -7304 50662 -7301
rect 50329 -7330 50470 -7304
rect 50277 -7363 50329 -7353
rect 50522 -7330 50662 -7304
rect 50470 -7366 50522 -7356
rect 50854 -7300 50906 -7293
rect 51046 -7298 51098 -7288
rect 50714 -7303 51046 -7300
rect 50714 -7330 50854 -7303
rect 50662 -7361 50714 -7351
rect 50906 -7330 51046 -7303
rect 50854 -7365 50906 -7355
rect 51238 -7299 51290 -7289
rect 51098 -7330 51238 -7300
rect 51046 -7360 51098 -7350
rect 51428 -7298 51480 -7288
rect 51290 -7330 51428 -7300
rect 51238 -7361 51290 -7351
rect 51622 -7300 51674 -7299
rect 51811 -7300 51863 -7297
rect 52000 -7300 52060 -6890
rect 52200 -7300 52252 -7298
rect 52390 -7300 52450 -6890
rect 52582 -7300 52634 -7298
rect 52774 -7300 52826 -7291
rect 52960 -7300 53020 -6890
rect 53159 -7300 53211 -7292
rect 53350 -7300 53410 -6890
rect 53542 -7300 53594 -7290
rect 53730 -7300 53790 -6890
rect 54120 -7287 54180 -6890
rect 53927 -7300 53979 -7291
rect 54119 -7297 54180 -7287
rect 54510 -7291 54570 -6890
rect 54890 -7290 54950 -6890
rect 55260 -7288 55320 -6890
rect 51480 -7301 53351 -7300
rect 51480 -7307 52774 -7301
rect 51480 -7309 51811 -7307
rect 51480 -7330 51622 -7309
rect 51428 -7360 51480 -7350
rect 51674 -7330 51811 -7309
rect 51622 -7371 51674 -7361
rect 51863 -7330 52001 -7307
rect 51811 -7369 51863 -7359
rect 52053 -7308 52392 -7307
rect 52053 -7330 52200 -7308
rect 52001 -7369 52053 -7359
rect 52252 -7330 52392 -7308
rect 52200 -7370 52252 -7360
rect 52444 -7308 52774 -7307
rect 52444 -7330 52582 -7308
rect 52392 -7369 52444 -7359
rect 52634 -7330 52774 -7308
rect 52582 -7370 52634 -7360
rect 52826 -7302 53351 -7301
rect 52826 -7303 53159 -7302
rect 52826 -7330 52966 -7303
rect 52774 -7363 52826 -7353
rect 53018 -7330 53159 -7303
rect 52966 -7365 53018 -7355
rect 53211 -7330 53351 -7302
rect 53159 -7364 53211 -7354
rect 53403 -7330 53542 -7300
rect 53351 -7362 53403 -7352
rect 53594 -7301 54119 -7300
rect 53594 -7305 53927 -7301
rect 53594 -7330 53736 -7305
rect 53542 -7362 53594 -7352
rect 53788 -7330 53927 -7305
rect 53736 -7367 53788 -7357
rect 53979 -7330 54119 -7301
rect 53927 -7363 53979 -7353
rect 54171 -7300 54180 -7297
rect 54312 -7300 54364 -7291
rect 54504 -7300 54570 -7291
rect 54697 -7300 54749 -7292
rect 54889 -7300 54950 -7290
rect 55080 -7299 55132 -7289
rect 54171 -7301 54889 -7300
rect 54171 -7330 54312 -7301
rect 54119 -7359 54171 -7349
rect 54364 -7330 54504 -7301
rect 54312 -7363 54364 -7353
rect 54556 -7302 54889 -7301
rect 54556 -7330 54697 -7302
rect 54504 -7363 54556 -7353
rect 54749 -7330 54889 -7302
rect 54697 -7364 54749 -7354
rect 54941 -7330 55080 -7300
rect 54889 -7362 54941 -7352
rect 55260 -7298 55323 -7288
rect 55260 -7300 55271 -7298
rect 55132 -7330 55271 -7300
rect 55080 -7361 55132 -7351
rect 55464 -7298 55516 -7288
rect 55323 -7330 55464 -7300
rect 55271 -7360 55323 -7350
rect 55650 -7300 55710 -6890
rect 55846 -7300 55898 -7298
rect 56030 -7300 56090 -6890
rect 56410 -7300 56470 -6890
rect 56810 -7300 56870 -6890
rect 57180 -7296 57240 -6890
rect 56997 -7300 57049 -7298
rect 57180 -7300 57243 -7296
rect 57384 -7300 57436 -7297
rect 57570 -7300 57630 -6890
rect 57960 -7298 58020 -6890
rect 57766 -7300 57818 -7298
rect 57959 -7300 58020 -7298
rect 58151 -7300 58203 -7298
rect 58340 -7300 58400 -6890
rect 58730 -7297 58790 -6890
rect 58535 -7300 58587 -7298
rect 58726 -7300 58790 -7297
rect 58921 -7300 58973 -7298
rect 59110 -7300 59170 -6890
rect 59303 -7300 59355 -7298
rect 59490 -7300 59550 -6890
rect 59880 -7298 59940 -6890
rect 59686 -7300 59738 -7298
rect 59878 -7300 59940 -7298
rect 60071 -7300 60123 -7298
rect 60260 -7300 60320 -6890
rect 60454 -7300 60506 -7298
rect 60640 -7300 60700 -6890
rect 60838 -7300 60890 -7298
rect 61030 -7300 61090 -6890
rect 61420 -7297 61480 -6890
rect 61222 -7300 61274 -7299
rect 61415 -7300 61480 -7297
rect 61605 -7300 61657 -7297
rect 61800 -7299 61860 -6890
rect 61798 -7300 61860 -7299
rect 61990 -7300 62042 -7298
rect 62180 -7300 62240 -6890
rect 62374 -7300 62426 -7297
rect 62570 -7298 62630 -6890
rect 62950 -7298 63010 -6890
rect 62566 -7300 62630 -7298
rect 62757 -7300 62809 -7298
rect 62949 -7300 63010 -7298
rect 63143 -7300 63195 -7297
rect 63340 -7298 63400 -6890
rect 63335 -7300 63400 -7298
rect 63525 -7300 63577 -7299
rect 63720 -7300 63780 -6890
rect 66912 -6912 66964 -6902
rect 63909 -7300 63961 -7298
rect 64102 -7300 64154 -7297
rect 64295 -7300 64347 -7298
rect 64486 -7300 64538 -7298
rect 64677 -7300 64729 -7298
rect 64870 -7300 64922 -7298
rect 65063 -7300 65115 -7298
rect 65254 -7300 65306 -7298
rect 65445 -7300 65497 -7297
rect 65636 -7300 65688 -7297
rect 65829 -7300 65881 -7298
rect 66023 -7300 66075 -7298
rect 66211 -7300 66263 -7299
rect 55516 -7306 66470 -7300
rect 55516 -7307 57191 -7306
rect 55516 -7330 55655 -7307
rect 55464 -7360 55516 -7350
rect 55707 -7308 57191 -7307
rect 55707 -7330 55846 -7308
rect 55655 -7369 55707 -7359
rect 55898 -7309 56997 -7308
rect 55898 -7330 56036 -7309
rect 55846 -7370 55898 -7360
rect 56088 -7311 56997 -7309
rect 56088 -7313 56808 -7311
rect 56088 -7330 56230 -7313
rect 56036 -7371 56088 -7361
rect 56282 -7314 56808 -7313
rect 56282 -7315 56616 -7314
rect 56282 -7330 56422 -7315
rect 56230 -7375 56282 -7365
rect 56474 -7330 56616 -7315
rect 56422 -7377 56474 -7367
rect 56668 -7330 56808 -7314
rect 56616 -7376 56668 -7366
rect 56860 -7330 56997 -7311
rect 56808 -7373 56860 -7363
rect 57049 -7330 57191 -7308
rect 56997 -7370 57049 -7360
rect 57243 -7307 66470 -7306
rect 57243 -7330 57384 -7307
rect 57191 -7368 57243 -7358
rect 57436 -7308 58726 -7307
rect 57436 -7330 57577 -7308
rect 57384 -7369 57436 -7359
rect 57629 -7330 57766 -7308
rect 57577 -7370 57629 -7360
rect 57818 -7330 57959 -7308
rect 57766 -7370 57818 -7360
rect 58011 -7330 58151 -7308
rect 57959 -7370 58011 -7360
rect 58203 -7330 58342 -7308
rect 58151 -7370 58203 -7360
rect 58394 -7330 58535 -7308
rect 58342 -7370 58394 -7360
rect 58587 -7330 58726 -7308
rect 58535 -7370 58587 -7360
rect 58778 -7308 61415 -7307
rect 58778 -7330 58921 -7308
rect 58726 -7369 58778 -7359
rect 58973 -7330 59110 -7308
rect 58921 -7370 58973 -7360
rect 59162 -7330 59303 -7308
rect 59110 -7370 59162 -7360
rect 59355 -7330 59495 -7308
rect 59303 -7370 59355 -7360
rect 59547 -7330 59686 -7308
rect 59495 -7370 59547 -7360
rect 59738 -7330 59878 -7308
rect 59686 -7370 59738 -7360
rect 59930 -7330 60071 -7308
rect 59878 -7370 59930 -7360
rect 60123 -7309 60454 -7308
rect 60123 -7330 60260 -7309
rect 60071 -7370 60123 -7360
rect 60312 -7330 60454 -7309
rect 60260 -7371 60312 -7361
rect 60506 -7330 60645 -7308
rect 60454 -7370 60506 -7360
rect 60697 -7330 60838 -7308
rect 60645 -7370 60697 -7360
rect 60890 -7330 61030 -7308
rect 60838 -7370 60890 -7360
rect 61082 -7309 61415 -7308
rect 61082 -7330 61222 -7309
rect 61030 -7370 61082 -7360
rect 61274 -7330 61415 -7309
rect 61222 -7371 61274 -7361
rect 61467 -7330 61605 -7307
rect 61415 -7369 61467 -7359
rect 61657 -7308 62183 -7307
rect 61657 -7309 61990 -7308
rect 61657 -7330 61798 -7309
rect 61605 -7369 61657 -7359
rect 61850 -7330 61990 -7309
rect 61798 -7371 61850 -7361
rect 62042 -7330 62183 -7308
rect 61990 -7370 62042 -7360
rect 62235 -7330 62374 -7307
rect 62183 -7369 62235 -7359
rect 62426 -7308 63143 -7307
rect 62426 -7330 62566 -7308
rect 62374 -7369 62426 -7359
rect 62618 -7330 62757 -7308
rect 62566 -7370 62618 -7360
rect 62809 -7330 62949 -7308
rect 62757 -7370 62809 -7360
rect 63001 -7330 63143 -7308
rect 62949 -7370 63001 -7360
rect 63195 -7308 64102 -7307
rect 63195 -7330 63335 -7308
rect 63143 -7369 63195 -7359
rect 63387 -7309 63909 -7308
rect 63387 -7330 63525 -7309
rect 63335 -7370 63387 -7360
rect 63577 -7310 63909 -7309
rect 63577 -7330 63716 -7310
rect 63525 -7371 63577 -7361
rect 63768 -7330 63909 -7310
rect 63716 -7372 63768 -7362
rect 63961 -7330 64102 -7308
rect 63909 -7370 63961 -7360
rect 64154 -7308 65445 -7307
rect 64154 -7330 64295 -7308
rect 64102 -7369 64154 -7359
rect 64347 -7330 64486 -7308
rect 64295 -7370 64347 -7360
rect 64538 -7330 64677 -7308
rect 64486 -7370 64538 -7360
rect 64729 -7330 64870 -7308
rect 64677 -7370 64729 -7360
rect 64922 -7330 65063 -7308
rect 64870 -7370 64922 -7360
rect 65115 -7330 65254 -7308
rect 65063 -7370 65115 -7360
rect 65306 -7330 65445 -7308
rect 65254 -7370 65306 -7360
rect 65497 -7330 65636 -7307
rect 65445 -7369 65497 -7359
rect 65688 -7308 66470 -7307
rect 65688 -7330 65829 -7308
rect 65636 -7369 65688 -7359
rect 65881 -7330 66023 -7308
rect 65829 -7370 65881 -7360
rect 66075 -7309 66470 -7308
rect 66075 -7330 66211 -7309
rect 66023 -7370 66075 -7360
rect 66263 -7317 66470 -7309
rect 66263 -7330 66405 -7317
rect 66211 -7371 66263 -7361
rect 66457 -7330 66470 -7317
rect 66405 -7379 66457 -7369
rect 49991 -7445 50043 -7435
rect 50182 -7447 50234 -7437
rect 50043 -7490 50182 -7460
rect 50043 -7497 50070 -7490
rect 49991 -7507 50070 -7497
rect 50000 -7654 50070 -7507
rect 50374 -7446 50426 -7436
rect 50234 -7490 50374 -7460
rect 50182 -7509 50234 -7499
rect 50566 -7449 50618 -7439
rect 50426 -7490 50566 -7460
rect 50374 -7508 50426 -7498
rect 50760 -7448 50812 -7438
rect 50618 -7490 50760 -7460
rect 50566 -7511 50618 -7501
rect 50950 -7448 51002 -7438
rect 50812 -7490 50950 -7460
rect 50760 -7510 50812 -7500
rect 51145 -7446 51197 -7436
rect 51002 -7490 51145 -7460
rect 50950 -7510 51002 -7500
rect 51336 -7445 51388 -7435
rect 51197 -7490 51336 -7460
rect 51145 -7508 51197 -7498
rect 51531 -7447 51583 -7437
rect 51388 -7490 51531 -7460
rect 51336 -7507 51388 -7497
rect 51721 -7447 51773 -7437
rect 51583 -7490 51721 -7460
rect 51531 -7509 51583 -7499
rect 51911 -7446 51963 -7436
rect 51773 -7490 51911 -7460
rect 51721 -7509 51773 -7499
rect 52104 -7445 52156 -7435
rect 51963 -7490 52104 -7460
rect 51911 -7508 51963 -7498
rect 52295 -7445 52347 -7435
rect 52156 -7490 52295 -7460
rect 52104 -7507 52156 -7497
rect 52491 -7447 52543 -7437
rect 52347 -7490 52491 -7460
rect 52295 -7507 52347 -7497
rect 52680 -7447 52732 -7437
rect 52543 -7490 52680 -7460
rect 52491 -7509 52543 -7499
rect 52874 -7447 52926 -7437
rect 52732 -7490 52874 -7460
rect 52680 -7509 52732 -7499
rect 53063 -7447 53115 -7437
rect 52926 -7490 53063 -7460
rect 52874 -7509 52926 -7499
rect 53255 -7448 53307 -7438
rect 53115 -7490 53255 -7460
rect 53063 -7509 53115 -7499
rect 53448 -7448 53500 -7438
rect 53307 -7490 53448 -7460
rect 53255 -7510 53307 -7500
rect 53639 -7448 53691 -7438
rect 53500 -7490 53639 -7460
rect 53448 -7510 53500 -7500
rect 53831 -7447 53883 -7437
rect 53691 -7490 53831 -7460
rect 53639 -7510 53691 -7500
rect 54023 -7448 54075 -7438
rect 53883 -7490 54023 -7460
rect 53831 -7509 53883 -7499
rect 54216 -7448 54268 -7438
rect 54075 -7490 54216 -7460
rect 54023 -7510 54075 -7500
rect 54407 -7448 54459 -7438
rect 54268 -7490 54407 -7460
rect 54216 -7510 54268 -7500
rect 54599 -7447 54651 -7437
rect 54459 -7490 54599 -7460
rect 54407 -7510 54459 -7500
rect 54792 -7448 54844 -7438
rect 54651 -7490 54792 -7460
rect 54599 -7509 54651 -7499
rect 54984 -7448 55036 -7438
rect 54844 -7490 54984 -7460
rect 54792 -7510 54844 -7500
rect 55175 -7448 55227 -7438
rect 55036 -7490 55175 -7460
rect 54984 -7510 55036 -7500
rect 55366 -7448 55418 -7438
rect 55227 -7490 55366 -7460
rect 55175 -7510 55227 -7500
rect 55558 -7448 55610 -7438
rect 55418 -7490 55558 -7460
rect 55366 -7510 55418 -7500
rect 55751 -7447 55803 -7437
rect 55610 -7490 55751 -7460
rect 55558 -7510 55610 -7500
rect 55942 -7447 55994 -7437
rect 55803 -7490 55942 -7460
rect 55751 -7509 55803 -7499
rect 56136 -7448 56188 -7438
rect 55994 -7490 56136 -7460
rect 55942 -7509 55994 -7499
rect 56328 -7448 56380 -7438
rect 56188 -7490 56328 -7460
rect 56136 -7510 56188 -7500
rect 56520 -7448 56572 -7438
rect 56380 -7490 56520 -7460
rect 56328 -7510 56380 -7500
rect 56712 -7448 56764 -7438
rect 56572 -7490 56712 -7460
rect 56520 -7510 56572 -7500
rect 56904 -7448 56956 -7438
rect 56764 -7490 56904 -7460
rect 56712 -7510 56764 -7500
rect 57096 -7448 57148 -7438
rect 56956 -7490 57096 -7460
rect 56904 -7510 56956 -7500
rect 57288 -7448 57340 -7438
rect 57148 -7490 57288 -7460
rect 57096 -7510 57148 -7500
rect 57479 -7448 57531 -7438
rect 57340 -7490 57479 -7460
rect 57288 -7510 57340 -7500
rect 57671 -7448 57723 -7438
rect 57531 -7490 57671 -7460
rect 57479 -7510 57531 -7500
rect 57864 -7448 57916 -7438
rect 57723 -7490 57864 -7460
rect 57671 -7510 57723 -7500
rect 58056 -7448 58108 -7438
rect 57916 -7490 58056 -7460
rect 57864 -7510 57916 -7500
rect 58248 -7448 58300 -7438
rect 58108 -7490 58248 -7460
rect 58056 -7510 58108 -7500
rect 58439 -7448 58491 -7438
rect 58300 -7490 58439 -7460
rect 58248 -7510 58300 -7500
rect 58631 -7448 58683 -7438
rect 58491 -7490 58631 -7460
rect 58439 -7510 58491 -7500
rect 58822 -7448 58874 -7438
rect 58683 -7490 58822 -7460
rect 58631 -7510 58683 -7500
rect 59013 -7448 59065 -7438
rect 58874 -7490 59013 -7460
rect 58822 -7510 58874 -7500
rect 59207 -7448 59259 -7438
rect 59065 -7490 59207 -7460
rect 59013 -7510 59065 -7500
rect 59399 -7448 59451 -7438
rect 59259 -7490 59399 -7460
rect 59207 -7510 59259 -7500
rect 59592 -7447 59644 -7437
rect 59451 -7490 59592 -7460
rect 59399 -7510 59451 -7500
rect 59783 -7448 59835 -7438
rect 59644 -7490 59783 -7460
rect 59592 -7509 59644 -7499
rect 59975 -7448 60027 -7438
rect 59835 -7490 59975 -7460
rect 59783 -7510 59835 -7500
rect 60168 -7448 60220 -7438
rect 60027 -7490 60168 -7460
rect 59975 -7510 60027 -7500
rect 60360 -7448 60412 -7438
rect 60220 -7490 60360 -7460
rect 60168 -7510 60220 -7500
rect 60553 -7447 60605 -7437
rect 60412 -7490 60553 -7460
rect 60360 -7510 60412 -7500
rect 60744 -7448 60796 -7438
rect 60605 -7490 60744 -7460
rect 60553 -7509 60605 -7499
rect 60936 -7448 60988 -7438
rect 60796 -7490 60936 -7460
rect 60744 -7510 60796 -7500
rect 61127 -7448 61179 -7438
rect 60988 -7490 61127 -7460
rect 60936 -7510 60988 -7500
rect 61319 -7448 61371 -7438
rect 61179 -7490 61319 -7460
rect 61127 -7510 61179 -7500
rect 61511 -7448 61563 -7438
rect 61371 -7490 61511 -7460
rect 61319 -7510 61371 -7500
rect 61704 -7448 61756 -7438
rect 61563 -7490 61704 -7460
rect 61511 -7510 61563 -7500
rect 61895 -7448 61947 -7438
rect 61756 -7490 61895 -7460
rect 61704 -7510 61756 -7500
rect 62087 -7448 62139 -7438
rect 61947 -7490 62087 -7460
rect 61895 -7510 61947 -7500
rect 62279 -7447 62331 -7437
rect 62139 -7490 62279 -7460
rect 62087 -7510 62139 -7500
rect 62471 -7448 62523 -7438
rect 62331 -7490 62471 -7460
rect 62279 -7509 62331 -7499
rect 62661 -7448 62713 -7438
rect 62523 -7490 62661 -7460
rect 62471 -7510 62523 -7500
rect 62855 -7448 62907 -7438
rect 62713 -7490 62855 -7460
rect 62661 -7510 62713 -7500
rect 63047 -7447 63099 -7437
rect 62907 -7490 63047 -7460
rect 62855 -7510 62907 -7500
rect 63238 -7448 63290 -7438
rect 63099 -7490 63238 -7460
rect 63047 -7509 63099 -7499
rect 63431 -7448 63483 -7438
rect 63290 -7490 63431 -7460
rect 63238 -7510 63290 -7500
rect 63622 -7447 63674 -7437
rect 63483 -7490 63622 -7460
rect 63431 -7510 63483 -7500
rect 63814 -7448 63866 -7438
rect 63674 -7490 63814 -7460
rect 63622 -7509 63674 -7499
rect 64005 -7448 64057 -7438
rect 63866 -7490 64005 -7460
rect 63814 -7510 63866 -7500
rect 64199 -7447 64251 -7437
rect 64057 -7490 64199 -7460
rect 64005 -7510 64057 -7500
rect 64390 -7448 64442 -7438
rect 64251 -7490 64390 -7460
rect 64199 -7509 64251 -7499
rect 64582 -7448 64634 -7438
rect 64442 -7490 64582 -7460
rect 64390 -7510 64442 -7500
rect 64774 -7448 64826 -7438
rect 64634 -7490 64774 -7460
rect 64582 -7510 64634 -7500
rect 64966 -7448 65018 -7438
rect 64826 -7490 64966 -7460
rect 64774 -7510 64826 -7500
rect 65159 -7448 65211 -7438
rect 65018 -7490 65159 -7460
rect 64966 -7510 65018 -7500
rect 65350 -7448 65402 -7438
rect 65211 -7490 65350 -7460
rect 65159 -7510 65211 -7500
rect 65543 -7447 65595 -7437
rect 65402 -7490 65543 -7460
rect 65350 -7510 65402 -7500
rect 65734 -7448 65786 -7438
rect 65595 -7490 65734 -7460
rect 65543 -7509 65595 -7499
rect 65927 -7448 65979 -7438
rect 65786 -7490 65927 -7460
rect 65734 -7510 65786 -7500
rect 66118 -7448 66170 -7438
rect 65979 -7490 66118 -7460
rect 65927 -7510 65979 -7500
rect 66309 -7446 66361 -7436
rect 66170 -7490 66309 -7460
rect 66118 -7510 66170 -7500
rect 66504 -7448 66556 -7438
rect 66361 -7490 66504 -7460
rect 66309 -7508 66361 -7498
rect 66440 -7500 66504 -7490
rect 66440 -7510 66556 -7500
rect 66440 -7654 66510 -7510
rect 49940 -7664 66588 -7654
rect 47224 -7808 47652 -7752
rect 48274 -7706 48446 -7696
rect 48274 -7774 48446 -7764
rect 49940 -7766 66588 -7756
rect 68120 -7710 68292 -7700
rect 68120 -7778 68292 -7768
rect 68894 -7756 68924 -6672
rect 69290 -7756 69326 -6672
rect 68894 -7806 69326 -7756
rect 68584 -7808 69326 -7806
rect 47224 -8196 69326 -7808
rect 47482 -8198 69326 -8196
<< via2 >>
rect 48274 -7764 48432 -7706
rect 49940 -7756 66574 -7664
rect 68120 -7768 68278 -7710
<< metal3 >>
rect 49104 -6370 49384 -6366
rect 52300 -6370 52394 -6366
rect 55614 -6370 55894 -6366
rect 62104 -6370 62384 -6366
rect 64654 -6370 64934 -6366
rect 67454 -6370 67734 -6366
rect 46324 -6434 51998 -6370
rect 52300 -6388 57790 -6370
rect 57908 -6388 58126 -6370
rect 52300 -6398 58126 -6388
rect 58606 -6398 69966 -6370
rect 52300 -6434 69966 -6398
rect 46324 -6648 69966 -6434
rect 49104 -7510 49384 -6648
rect 52114 -7510 52394 -6648
rect 55614 -7510 55894 -6648
rect 62104 -7510 62384 -6648
rect 64654 -7510 64934 -6648
rect 67454 -7510 67734 -6648
rect 46350 -7664 69992 -7510
rect 46350 -7706 49940 -7664
rect 46350 -7764 48274 -7706
rect 48432 -7756 49940 -7706
rect 66574 -7710 69992 -7664
rect 66574 -7756 68120 -7710
rect 48432 -7764 68120 -7756
rect 46350 -7768 68120 -7764
rect 68278 -7768 69992 -7710
rect 46350 -7788 69992 -7768
use sky130_fd_pr__nfet_01v8_lvt_FKGFGD  XM20
timestamp 1662412052
transform 1 0 54905 0 1 -6780
box -3095 -310 3095 310
use sky130_fd_pr__nfet_01v8_lvt_FKGFGD  XM23
timestamp 1662412052
transform 1 0 61095 0 1 -6780
box -3095 -310 3095 310
use sky130_fd_pr__nfet_01v8_lvt_G3ZQK6  XM25
timestamp 1662412052
transform 1 0 58273 0 1 -7398
box -8423 -310 8423 310
use sky130_fd_pr__res_xhigh_po_5p73_4C7XCD  XR19
timestamp 1662952458
transform 0 1 47715 -1 0 -7211
box -739 -657 739 657
use sky130_fd_pr__nfet_01v8_lvt_HFYJAZ  sky130_fd_pr__nfet_01v8_lvt_HFYJAZ_0
timestamp 1662983156
transform 1 0 49649 0 1 -7275
box -211 -447 211 447
use sky130_fd_pr__res_high_po_0p35_C28PVF  sky130_fd_pr__res_high_po_0p35_C28PVF_0
timestamp 1662983156
transform 1 0 48973 0 1 -6540
box -201 -998 201 998
use sky130_fd_pr__res_high_po_0p35_C28PVF  sky130_fd_pr__res_high_po_0p35_C28PVF_1
timestamp 1662983156
transform 1 0 67579 0 1 -6624
box -201 -998 201 998
use sky130_fd_pr__res_xhigh_po_5p73_4C7XCD  sky130_fd_pr__res_xhigh_po_5p73_4C7XCD_0
timestamp 1662952458
transform 0 1 68837 -1 0 -7211
box -739 -657 739 657
<< labels >>
rlabel metal2 47482 -8198 69326 -7808 0 vdd
rlabel metal3 46324 -6648 51998 -6370 0 vss
rlabel metal1 49672 -7584 49724 -6302 0 Iref
rlabel metal1 51874 -6950 51904 -6358 0 vout5p
rlabel metal1 64088 -6944 64118 -6352 0 vout5n
rlabel metal1 48934 -5718 49008 -5432 0 vin0p
rlabel metal1 67544 -5802 67616 -5516 0 vin0n
<< end >>
