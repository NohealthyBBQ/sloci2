magic
tech sky130A
magscale 1 2
timestamp 1662761135
<< nwell >>
rect -683 -1191 683 1191
<< pmoslvt >>
rect -487 772 -287 972
rect -229 772 -29 972
rect 29 772 229 972
rect 287 772 487 972
rect -487 336 -287 536
rect -229 336 -29 536
rect 29 336 229 536
rect 287 336 487 536
rect -487 -100 -287 100
rect -229 -100 -29 100
rect 29 -100 229 100
rect 287 -100 487 100
rect -487 -536 -287 -336
rect -229 -536 -29 -336
rect 29 -536 229 -336
rect 287 -536 487 -336
rect -487 -972 -287 -772
rect -229 -972 -29 -772
rect 29 -972 229 -772
rect 287 -972 487 -772
<< pdiff >>
rect -545 960 -487 972
rect -545 784 -533 960
rect -499 784 -487 960
rect -545 772 -487 784
rect -287 960 -229 972
rect -287 784 -275 960
rect -241 784 -229 960
rect -287 772 -229 784
rect -29 960 29 972
rect -29 784 -17 960
rect 17 784 29 960
rect -29 772 29 784
rect 229 960 287 972
rect 229 784 241 960
rect 275 784 287 960
rect 229 772 287 784
rect 487 960 545 972
rect 487 784 499 960
rect 533 784 545 960
rect 487 772 545 784
rect -545 524 -487 536
rect -545 348 -533 524
rect -499 348 -487 524
rect -545 336 -487 348
rect -287 524 -229 536
rect -287 348 -275 524
rect -241 348 -229 524
rect -287 336 -229 348
rect -29 524 29 536
rect -29 348 -17 524
rect 17 348 29 524
rect -29 336 29 348
rect 229 524 287 536
rect 229 348 241 524
rect 275 348 287 524
rect 229 336 287 348
rect 487 524 545 536
rect 487 348 499 524
rect 533 348 545 524
rect 487 336 545 348
rect -545 88 -487 100
rect -545 -88 -533 88
rect -499 -88 -487 88
rect -545 -100 -487 -88
rect -287 88 -229 100
rect -287 -88 -275 88
rect -241 -88 -229 88
rect -287 -100 -229 -88
rect -29 88 29 100
rect -29 -88 -17 88
rect 17 -88 29 88
rect -29 -100 29 -88
rect 229 88 287 100
rect 229 -88 241 88
rect 275 -88 287 88
rect 229 -100 287 -88
rect 487 88 545 100
rect 487 -88 499 88
rect 533 -88 545 88
rect 487 -100 545 -88
rect -545 -348 -487 -336
rect -545 -524 -533 -348
rect -499 -524 -487 -348
rect -545 -536 -487 -524
rect -287 -348 -229 -336
rect -287 -524 -275 -348
rect -241 -524 -229 -348
rect -287 -536 -229 -524
rect -29 -348 29 -336
rect -29 -524 -17 -348
rect 17 -524 29 -348
rect -29 -536 29 -524
rect 229 -348 287 -336
rect 229 -524 241 -348
rect 275 -524 287 -348
rect 229 -536 287 -524
rect 487 -348 545 -336
rect 487 -524 499 -348
rect 533 -524 545 -348
rect 487 -536 545 -524
rect -545 -784 -487 -772
rect -545 -960 -533 -784
rect -499 -960 -487 -784
rect -545 -972 -487 -960
rect -287 -784 -229 -772
rect -287 -960 -275 -784
rect -241 -960 -229 -784
rect -287 -972 -229 -960
rect -29 -784 29 -772
rect -29 -960 -17 -784
rect 17 -960 29 -784
rect -29 -972 29 -960
rect 229 -784 287 -772
rect 229 -960 241 -784
rect 275 -960 287 -784
rect 229 -972 287 -960
rect 487 -784 545 -772
rect 487 -960 499 -784
rect 533 -960 545 -784
rect 487 -972 545 -960
<< pdiffc >>
rect -533 784 -499 960
rect -275 784 -241 960
rect -17 784 17 960
rect 241 784 275 960
rect 499 784 533 960
rect -533 348 -499 524
rect -275 348 -241 524
rect -17 348 17 524
rect 241 348 275 524
rect 499 348 533 524
rect -533 -88 -499 88
rect -275 -88 -241 88
rect -17 -88 17 88
rect 241 -88 275 88
rect 499 -88 533 88
rect -533 -524 -499 -348
rect -275 -524 -241 -348
rect -17 -524 17 -348
rect 241 -524 275 -348
rect 499 -524 533 -348
rect -533 -960 -499 -784
rect -275 -960 -241 -784
rect -17 -960 17 -784
rect 241 -960 275 -784
rect 499 -960 533 -784
<< nsubdiff >>
rect -647 1121 -551 1155
rect 551 1121 647 1155
rect -647 1059 -613 1121
rect 613 1059 647 1121
rect -647 -1121 -613 -1059
rect 613 -1121 647 -1059
rect -647 -1155 -551 -1121
rect 551 -1155 647 -1121
<< nsubdiffcont >>
rect -551 1121 551 1155
rect -647 -1059 -613 1059
rect 613 -1059 647 1059
rect -551 -1155 551 -1121
<< poly >>
rect -487 1053 -287 1069
rect -487 1019 -471 1053
rect -303 1019 -287 1053
rect -487 972 -287 1019
rect -229 1053 -29 1069
rect -229 1019 -213 1053
rect -45 1019 -29 1053
rect -229 972 -29 1019
rect 29 1053 229 1069
rect 29 1019 45 1053
rect 213 1019 229 1053
rect 29 972 229 1019
rect 287 1053 487 1069
rect 287 1019 303 1053
rect 471 1019 487 1053
rect 287 972 487 1019
rect -487 725 -287 772
rect -487 691 -471 725
rect -303 691 -287 725
rect -487 675 -287 691
rect -229 725 -29 772
rect -229 691 -213 725
rect -45 691 -29 725
rect -229 675 -29 691
rect 29 725 229 772
rect 29 691 45 725
rect 213 691 229 725
rect 29 675 229 691
rect 287 725 487 772
rect 287 691 303 725
rect 471 691 487 725
rect 287 675 487 691
rect -487 617 -287 633
rect -487 583 -471 617
rect -303 583 -287 617
rect -487 536 -287 583
rect -229 617 -29 633
rect -229 583 -213 617
rect -45 583 -29 617
rect -229 536 -29 583
rect 29 617 229 633
rect 29 583 45 617
rect 213 583 229 617
rect 29 536 229 583
rect 287 617 487 633
rect 287 583 303 617
rect 471 583 487 617
rect 287 536 487 583
rect -487 289 -287 336
rect -487 255 -471 289
rect -303 255 -287 289
rect -487 239 -287 255
rect -229 289 -29 336
rect -229 255 -213 289
rect -45 255 -29 289
rect -229 239 -29 255
rect 29 289 229 336
rect 29 255 45 289
rect 213 255 229 289
rect 29 239 229 255
rect 287 289 487 336
rect 287 255 303 289
rect 471 255 487 289
rect 287 239 487 255
rect -487 181 -287 197
rect -487 147 -471 181
rect -303 147 -287 181
rect -487 100 -287 147
rect -229 181 -29 197
rect -229 147 -213 181
rect -45 147 -29 181
rect -229 100 -29 147
rect 29 181 229 197
rect 29 147 45 181
rect 213 147 229 181
rect 29 100 229 147
rect 287 181 487 197
rect 287 147 303 181
rect 471 147 487 181
rect 287 100 487 147
rect -487 -147 -287 -100
rect -487 -181 -471 -147
rect -303 -181 -287 -147
rect -487 -197 -287 -181
rect -229 -147 -29 -100
rect -229 -181 -213 -147
rect -45 -181 -29 -147
rect -229 -197 -29 -181
rect 29 -147 229 -100
rect 29 -181 45 -147
rect 213 -181 229 -147
rect 29 -197 229 -181
rect 287 -147 487 -100
rect 287 -181 303 -147
rect 471 -181 487 -147
rect 287 -197 487 -181
rect -487 -255 -287 -239
rect -487 -289 -471 -255
rect -303 -289 -287 -255
rect -487 -336 -287 -289
rect -229 -255 -29 -239
rect -229 -289 -213 -255
rect -45 -289 -29 -255
rect -229 -336 -29 -289
rect 29 -255 229 -239
rect 29 -289 45 -255
rect 213 -289 229 -255
rect 29 -336 229 -289
rect 287 -255 487 -239
rect 287 -289 303 -255
rect 471 -289 487 -255
rect 287 -336 487 -289
rect -487 -583 -287 -536
rect -487 -617 -471 -583
rect -303 -617 -287 -583
rect -487 -633 -287 -617
rect -229 -583 -29 -536
rect -229 -617 -213 -583
rect -45 -617 -29 -583
rect -229 -633 -29 -617
rect 29 -583 229 -536
rect 29 -617 45 -583
rect 213 -617 229 -583
rect 29 -633 229 -617
rect 287 -583 487 -536
rect 287 -617 303 -583
rect 471 -617 487 -583
rect 287 -633 487 -617
rect -487 -691 -287 -675
rect -487 -725 -471 -691
rect -303 -725 -287 -691
rect -487 -772 -287 -725
rect -229 -691 -29 -675
rect -229 -725 -213 -691
rect -45 -725 -29 -691
rect -229 -772 -29 -725
rect 29 -691 229 -675
rect 29 -725 45 -691
rect 213 -725 229 -691
rect 29 -772 229 -725
rect 287 -691 487 -675
rect 287 -725 303 -691
rect 471 -725 487 -691
rect 287 -772 487 -725
rect -487 -1019 -287 -972
rect -487 -1053 -471 -1019
rect -303 -1053 -287 -1019
rect -487 -1069 -287 -1053
rect -229 -1019 -29 -972
rect -229 -1053 -213 -1019
rect -45 -1053 -29 -1019
rect -229 -1069 -29 -1053
rect 29 -1019 229 -972
rect 29 -1053 45 -1019
rect 213 -1053 229 -1019
rect 29 -1069 229 -1053
rect 287 -1019 487 -972
rect 287 -1053 303 -1019
rect 471 -1053 487 -1019
rect 287 -1069 487 -1053
<< polycont >>
rect -471 1019 -303 1053
rect -213 1019 -45 1053
rect 45 1019 213 1053
rect 303 1019 471 1053
rect -471 691 -303 725
rect -213 691 -45 725
rect 45 691 213 725
rect 303 691 471 725
rect -471 583 -303 617
rect -213 583 -45 617
rect 45 583 213 617
rect 303 583 471 617
rect -471 255 -303 289
rect -213 255 -45 289
rect 45 255 213 289
rect 303 255 471 289
rect -471 147 -303 181
rect -213 147 -45 181
rect 45 147 213 181
rect 303 147 471 181
rect -471 -181 -303 -147
rect -213 -181 -45 -147
rect 45 -181 213 -147
rect 303 -181 471 -147
rect -471 -289 -303 -255
rect -213 -289 -45 -255
rect 45 -289 213 -255
rect 303 -289 471 -255
rect -471 -617 -303 -583
rect -213 -617 -45 -583
rect 45 -617 213 -583
rect 303 -617 471 -583
rect -471 -725 -303 -691
rect -213 -725 -45 -691
rect 45 -725 213 -691
rect 303 -725 471 -691
rect -471 -1053 -303 -1019
rect -213 -1053 -45 -1019
rect 45 -1053 213 -1019
rect 303 -1053 471 -1019
<< locali >>
rect -647 1121 -551 1155
rect 551 1121 647 1155
rect -647 1059 -613 1121
rect 613 1059 647 1121
rect -487 1019 -471 1053
rect -303 1019 -287 1053
rect -229 1019 -213 1053
rect -45 1019 -29 1053
rect 29 1019 45 1053
rect 213 1019 229 1053
rect 287 1019 303 1053
rect 471 1019 487 1053
rect -533 960 -499 976
rect -533 768 -499 784
rect -275 960 -241 976
rect -275 768 -241 784
rect -17 960 17 976
rect -17 768 17 784
rect 241 960 275 976
rect 241 768 275 784
rect 499 960 533 976
rect 499 768 533 784
rect -487 691 -471 725
rect -303 691 -287 725
rect -229 691 -213 725
rect -45 691 -29 725
rect 29 691 45 725
rect 213 691 229 725
rect 287 691 303 725
rect 471 691 487 725
rect -487 583 -471 617
rect -303 583 -287 617
rect -229 583 -213 617
rect -45 583 -29 617
rect 29 583 45 617
rect 213 583 229 617
rect 287 583 303 617
rect 471 583 487 617
rect -533 524 -499 540
rect -533 332 -499 348
rect -275 524 -241 540
rect -275 332 -241 348
rect -17 524 17 540
rect -17 332 17 348
rect 241 524 275 540
rect 241 332 275 348
rect 499 524 533 540
rect 499 332 533 348
rect -487 255 -471 289
rect -303 255 -287 289
rect -229 255 -213 289
rect -45 255 -29 289
rect 29 255 45 289
rect 213 255 229 289
rect 287 255 303 289
rect 471 255 487 289
rect -487 147 -471 181
rect -303 147 -287 181
rect -229 147 -213 181
rect -45 147 -29 181
rect 29 147 45 181
rect 213 147 229 181
rect 287 147 303 181
rect 471 147 487 181
rect -533 88 -499 104
rect -533 -104 -499 -88
rect -275 88 -241 104
rect -275 -104 -241 -88
rect -17 88 17 104
rect -17 -104 17 -88
rect 241 88 275 104
rect 241 -104 275 -88
rect 499 88 533 104
rect 499 -104 533 -88
rect -487 -181 -471 -147
rect -303 -181 -287 -147
rect -229 -181 -213 -147
rect -45 -181 -29 -147
rect 29 -181 45 -147
rect 213 -181 229 -147
rect 287 -181 303 -147
rect 471 -181 487 -147
rect -487 -289 -471 -255
rect -303 -289 -287 -255
rect -229 -289 -213 -255
rect -45 -289 -29 -255
rect 29 -289 45 -255
rect 213 -289 229 -255
rect 287 -289 303 -255
rect 471 -289 487 -255
rect -533 -348 -499 -332
rect -533 -540 -499 -524
rect -275 -348 -241 -332
rect -275 -540 -241 -524
rect -17 -348 17 -332
rect -17 -540 17 -524
rect 241 -348 275 -332
rect 241 -540 275 -524
rect 499 -348 533 -332
rect 499 -540 533 -524
rect -487 -617 -471 -583
rect -303 -617 -287 -583
rect -229 -617 -213 -583
rect -45 -617 -29 -583
rect 29 -617 45 -583
rect 213 -617 229 -583
rect 287 -617 303 -583
rect 471 -617 487 -583
rect -487 -725 -471 -691
rect -303 -725 -287 -691
rect -229 -725 -213 -691
rect -45 -725 -29 -691
rect 29 -725 45 -691
rect 213 -725 229 -691
rect 287 -725 303 -691
rect 471 -725 487 -691
rect -533 -784 -499 -768
rect -533 -976 -499 -960
rect -275 -784 -241 -768
rect -275 -976 -241 -960
rect -17 -784 17 -768
rect -17 -976 17 -960
rect 241 -784 275 -768
rect 241 -976 275 -960
rect 499 -784 533 -768
rect 499 -976 533 -960
rect -487 -1053 -471 -1019
rect -303 -1053 -287 -1019
rect -229 -1053 -213 -1019
rect -45 -1053 -29 -1019
rect 29 -1053 45 -1019
rect 213 -1053 229 -1019
rect 287 -1053 303 -1019
rect 471 -1053 487 -1019
rect -647 -1121 -613 -1059
rect 613 -1121 647 -1059
rect -647 -1155 -551 -1121
rect 551 -1155 647 -1121
<< viali >>
rect -471 1019 -303 1053
rect -213 1019 -45 1053
rect 45 1019 213 1053
rect 303 1019 471 1053
rect -533 784 -499 960
rect -275 784 -241 960
rect -17 784 17 960
rect 241 784 275 960
rect 499 784 533 960
rect -471 691 -303 725
rect -213 691 -45 725
rect 45 691 213 725
rect 303 691 471 725
rect -471 583 -303 617
rect -213 583 -45 617
rect 45 583 213 617
rect 303 583 471 617
rect -533 348 -499 524
rect -275 348 -241 524
rect -17 348 17 524
rect 241 348 275 524
rect 499 348 533 524
rect -471 255 -303 289
rect -213 255 -45 289
rect 45 255 213 289
rect 303 255 471 289
rect -471 147 -303 181
rect -213 147 -45 181
rect 45 147 213 181
rect 303 147 471 181
rect -533 -88 -499 88
rect -275 -88 -241 88
rect -17 -88 17 88
rect 241 -88 275 88
rect 499 -88 533 88
rect -471 -181 -303 -147
rect -213 -181 -45 -147
rect 45 -181 213 -147
rect 303 -181 471 -147
rect -471 -289 -303 -255
rect -213 -289 -45 -255
rect 45 -289 213 -255
rect 303 -289 471 -255
rect -533 -524 -499 -348
rect -275 -524 -241 -348
rect -17 -524 17 -348
rect 241 -524 275 -348
rect 499 -524 533 -348
rect -471 -617 -303 -583
rect -213 -617 -45 -583
rect 45 -617 213 -583
rect 303 -617 471 -583
rect -471 -725 -303 -691
rect -213 -725 -45 -691
rect 45 -725 213 -691
rect 303 -725 471 -691
rect -533 -960 -499 -784
rect -275 -960 -241 -784
rect -17 -960 17 -784
rect 241 -960 275 -784
rect 499 -960 533 -784
rect -471 -1053 -303 -1019
rect -213 -1053 -45 -1019
rect 45 -1053 213 -1019
rect 303 -1053 471 -1019
<< metal1 >>
rect -483 1053 -291 1059
rect -483 1019 -471 1053
rect -303 1019 -291 1053
rect -483 1013 -291 1019
rect -225 1053 -33 1059
rect -225 1019 -213 1053
rect -45 1019 -33 1053
rect -225 1013 -33 1019
rect 33 1053 225 1059
rect 33 1019 45 1053
rect 213 1019 225 1053
rect 33 1013 225 1019
rect 291 1053 483 1059
rect 291 1019 303 1053
rect 471 1019 483 1053
rect 291 1013 483 1019
rect -539 960 -493 972
rect -539 784 -533 960
rect -499 784 -493 960
rect -539 772 -493 784
rect -281 960 -235 972
rect -281 784 -275 960
rect -241 784 -235 960
rect -281 772 -235 784
rect -23 960 23 972
rect -23 784 -17 960
rect 17 784 23 960
rect -23 772 23 784
rect 235 960 281 972
rect 235 784 241 960
rect 275 784 281 960
rect 235 772 281 784
rect 493 960 539 972
rect 493 784 499 960
rect 533 784 539 960
rect 493 772 539 784
rect -483 725 -291 731
rect -483 691 -471 725
rect -303 691 -291 725
rect -483 685 -291 691
rect -225 725 -33 731
rect -225 691 -213 725
rect -45 691 -33 725
rect -225 685 -33 691
rect 33 725 225 731
rect 33 691 45 725
rect 213 691 225 725
rect 33 685 225 691
rect 291 725 483 731
rect 291 691 303 725
rect 471 691 483 725
rect 291 685 483 691
rect -483 617 -291 623
rect -483 583 -471 617
rect -303 583 -291 617
rect -483 577 -291 583
rect -225 617 -33 623
rect -225 583 -213 617
rect -45 583 -33 617
rect -225 577 -33 583
rect 33 617 225 623
rect 33 583 45 617
rect 213 583 225 617
rect 33 577 225 583
rect 291 617 483 623
rect 291 583 303 617
rect 471 583 483 617
rect 291 577 483 583
rect -539 524 -493 536
rect -539 348 -533 524
rect -499 348 -493 524
rect -539 336 -493 348
rect -281 524 -235 536
rect -281 348 -275 524
rect -241 348 -235 524
rect -281 336 -235 348
rect -23 524 23 536
rect -23 348 -17 524
rect 17 348 23 524
rect -23 336 23 348
rect 235 524 281 536
rect 235 348 241 524
rect 275 348 281 524
rect 235 336 281 348
rect 493 524 539 536
rect 493 348 499 524
rect 533 348 539 524
rect 493 336 539 348
rect -483 289 -291 295
rect -483 255 -471 289
rect -303 255 -291 289
rect -483 249 -291 255
rect -225 289 -33 295
rect -225 255 -213 289
rect -45 255 -33 289
rect -225 249 -33 255
rect 33 289 225 295
rect 33 255 45 289
rect 213 255 225 289
rect 33 249 225 255
rect 291 289 483 295
rect 291 255 303 289
rect 471 255 483 289
rect 291 249 483 255
rect -483 181 -291 187
rect -483 147 -471 181
rect -303 147 -291 181
rect -483 141 -291 147
rect -225 181 -33 187
rect -225 147 -213 181
rect -45 147 -33 181
rect -225 141 -33 147
rect 33 181 225 187
rect 33 147 45 181
rect 213 147 225 181
rect 33 141 225 147
rect 291 181 483 187
rect 291 147 303 181
rect 471 147 483 181
rect 291 141 483 147
rect -539 88 -493 100
rect -539 -88 -533 88
rect -499 -88 -493 88
rect -539 -100 -493 -88
rect -281 88 -235 100
rect -281 -88 -275 88
rect -241 -88 -235 88
rect -281 -100 -235 -88
rect -23 88 23 100
rect -23 -88 -17 88
rect 17 -88 23 88
rect -23 -100 23 -88
rect 235 88 281 100
rect 235 -88 241 88
rect 275 -88 281 88
rect 235 -100 281 -88
rect 493 88 539 100
rect 493 -88 499 88
rect 533 -88 539 88
rect 493 -100 539 -88
rect -483 -147 -291 -141
rect -483 -181 -471 -147
rect -303 -181 -291 -147
rect -483 -187 -291 -181
rect -225 -147 -33 -141
rect -225 -181 -213 -147
rect -45 -181 -33 -147
rect -225 -187 -33 -181
rect 33 -147 225 -141
rect 33 -181 45 -147
rect 213 -181 225 -147
rect 33 -187 225 -181
rect 291 -147 483 -141
rect 291 -181 303 -147
rect 471 -181 483 -147
rect 291 -187 483 -181
rect -483 -255 -291 -249
rect -483 -289 -471 -255
rect -303 -289 -291 -255
rect -483 -295 -291 -289
rect -225 -255 -33 -249
rect -225 -289 -213 -255
rect -45 -289 -33 -255
rect -225 -295 -33 -289
rect 33 -255 225 -249
rect 33 -289 45 -255
rect 213 -289 225 -255
rect 33 -295 225 -289
rect 291 -255 483 -249
rect 291 -289 303 -255
rect 471 -289 483 -255
rect 291 -295 483 -289
rect -539 -348 -493 -336
rect -539 -524 -533 -348
rect -499 -524 -493 -348
rect -539 -536 -493 -524
rect -281 -348 -235 -336
rect -281 -524 -275 -348
rect -241 -524 -235 -348
rect -281 -536 -235 -524
rect -23 -348 23 -336
rect -23 -524 -17 -348
rect 17 -524 23 -348
rect -23 -536 23 -524
rect 235 -348 281 -336
rect 235 -524 241 -348
rect 275 -524 281 -348
rect 235 -536 281 -524
rect 493 -348 539 -336
rect 493 -524 499 -348
rect 533 -524 539 -348
rect 493 -536 539 -524
rect -483 -583 -291 -577
rect -483 -617 -471 -583
rect -303 -617 -291 -583
rect -483 -623 -291 -617
rect -225 -583 -33 -577
rect -225 -617 -213 -583
rect -45 -617 -33 -583
rect -225 -623 -33 -617
rect 33 -583 225 -577
rect 33 -617 45 -583
rect 213 -617 225 -583
rect 33 -623 225 -617
rect 291 -583 483 -577
rect 291 -617 303 -583
rect 471 -617 483 -583
rect 291 -623 483 -617
rect -483 -691 -291 -685
rect -483 -725 -471 -691
rect -303 -725 -291 -691
rect -483 -731 -291 -725
rect -225 -691 -33 -685
rect -225 -725 -213 -691
rect -45 -725 -33 -691
rect -225 -731 -33 -725
rect 33 -691 225 -685
rect 33 -725 45 -691
rect 213 -725 225 -691
rect 33 -731 225 -725
rect 291 -691 483 -685
rect 291 -725 303 -691
rect 471 -725 483 -691
rect 291 -731 483 -725
rect -539 -784 -493 -772
rect -539 -960 -533 -784
rect -499 -960 -493 -784
rect -539 -972 -493 -960
rect -281 -784 -235 -772
rect -281 -960 -275 -784
rect -241 -960 -235 -784
rect -281 -972 -235 -960
rect -23 -784 23 -772
rect -23 -960 -17 -784
rect 17 -960 23 -784
rect -23 -972 23 -960
rect 235 -784 281 -772
rect 235 -960 241 -784
rect 275 -960 281 -784
rect 235 -972 281 -960
rect 493 -784 539 -772
rect 493 -960 499 -784
rect 533 -960 539 -784
rect 493 -972 539 -960
rect -483 -1019 -291 -1013
rect -483 -1053 -471 -1019
rect -303 -1053 -291 -1019
rect -483 -1059 -291 -1053
rect -225 -1019 -33 -1013
rect -225 -1053 -213 -1019
rect -45 -1053 -33 -1019
rect -225 -1059 -33 -1053
rect 33 -1019 225 -1013
rect 33 -1053 45 -1019
rect 213 -1053 225 -1019
rect 33 -1059 225 -1053
rect 291 -1019 483 -1013
rect 291 -1053 303 -1019
rect 471 -1053 483 -1019
rect 291 -1059 483 -1053
<< properties >>
string FIXED_BBOX -630 -1138 630 1138
string gencell sky130_fd_pr__pfet_01v8_lvt
string library sky130
string parameters w 1 l 1 m 5 nf 4 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.35 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
