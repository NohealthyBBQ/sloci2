magic
tech sky130A
magscale 1 2
timestamp 1672340817
<< metal1 >>
rect -960 3080 60 3100
rect -960 2980 -940 3080
rect -840 2980 60 3080
rect -960 2960 60 2980
rect 890 2660 900 2860
rect 1100 2660 1110 2860
rect -60 2160 100 2180
rect -60 2060 -40 2160
rect 60 2060 100 2160
rect -60 2040 100 2060
rect -300 1860 300 1900
rect -300 1740 -260 1860
rect -140 1740 300 1860
rect -300 1700 300 1740
rect 3380 -2380 3560 -2360
rect 3380 -2440 3480 -2380
rect 3540 -2440 3560 -2380
rect 3380 -2460 3560 -2440
rect 3260 -5220 3420 -4560
rect 3260 -5340 3280 -5220
rect 3400 -5340 3420 -5220
rect 3260 -5380 3420 -5340
rect -960 -24920 360 -24900
rect -960 -25020 -940 -24920
rect -840 -25020 360 -24920
rect -960 -25040 360 -25020
rect 1070 -25320 1080 -25120
rect 1360 -25320 1370 -25120
rect -580 -25840 300 -25820
rect -580 -25940 -560 -25840
rect -420 -25940 300 -25840
rect -580 -25960 300 -25940
rect -340 -26160 520 -26120
rect -340 -26340 -300 -26160
rect -160 -26340 520 -26160
rect -340 -26380 520 -26340
rect -960 -52520 220 -52500
rect -960 -52620 -940 -52520
rect -840 -52620 220 -52520
rect -960 -52640 220 -52620
rect -60 -53440 80 -53420
rect -60 -53540 -40 -53440
rect 60 -53540 80 -53440
rect -60 -53560 80 -53540
rect -340 -53780 320 -53740
rect -340 -53940 -300 -53780
rect -160 -53940 320 -53780
rect -340 -53980 320 -53940
<< via1 >>
rect -940 2980 -840 3080
rect 900 2660 1100 2860
rect -40 2060 60 2160
rect -260 1740 -140 1860
rect 3480 -2440 3540 -2380
rect 3280 -5340 3400 -5220
rect -940 -25020 -840 -24920
rect 1080 -25320 1360 -25120
rect -560 -25940 -420 -25840
rect -300 -26340 -160 -26160
rect -940 -52620 -840 -52520
rect -40 -53540 60 -53440
rect -300 -53940 -160 -53780
<< metal2 >>
rect -1100 3080 -700 3200
rect -1100 2980 -940 3080
rect -840 2980 -700 3080
rect -1100 -24920 -700 2980
rect 900 2860 1100 2870
rect 900 2650 1100 2660
rect -60 2160 80 2180
rect -60 2060 -40 2160
rect 60 2060 80 2160
rect -260 1860 -140 1870
rect -260 1730 -140 1740
rect -60 -1000 80 2060
rect -60 -1140 3560 -1000
rect 3460 -2380 3560 -1140
rect 3460 -2440 3480 -2380
rect 3540 -2440 3560 -2380
rect 3460 -2460 3560 -2440
rect 3340 -3440 3680 -3280
rect 3540 -5000 3680 -3440
rect -1100 -25020 -940 -24920
rect -840 -25020 -700 -24920
rect -1100 -52520 -700 -25020
rect -560 -5140 3680 -5000
rect -560 -25840 -420 -5140
rect -560 -25960 -420 -25940
rect -60 -5220 3420 -5200
rect -60 -5340 3280 -5220
rect 3400 -5340 3420 -5220
rect -60 -5360 3420 -5340
rect -300 -26160 -160 -26150
rect -300 -26350 -160 -26340
rect -1100 -52620 -940 -52520
rect -840 -52620 -700 -52520
rect -1100 -52700 -700 -52620
rect -60 -53440 80 -5360
rect 1080 -25120 1360 -25110
rect 1080 -25330 1360 -25320
rect -60 -53540 -40 -53440
rect 60 -53540 80 -53440
rect -60 -53560 80 -53540
rect -300 -53780 -160 -53770
rect -300 -53950 -160 -53940
<< via2 >>
rect 900 2660 1100 2860
rect -260 1740 -140 1860
rect -300 -26340 -160 -26160
rect 1080 -25320 1360 -25120
rect -300 -53940 -160 -53780
<< metal3 >>
rect 890 2860 1110 2865
rect 890 2660 900 2860
rect 1100 2660 1110 2860
rect 890 2655 1110 2660
rect -380 1860 -100 2440
rect -380 1740 -260 1860
rect -140 1740 -100 1860
rect -380 -26160 -100 1740
rect 1070 -25120 1370 -25115
rect 1070 -25320 1080 -25120
rect 1360 -25320 1370 -25120
rect 1070 -25325 1370 -25320
rect -380 -26340 -300 -26160
rect -160 -26340 -100 -26160
rect -380 -53780 -100 -26340
rect -380 -53940 -300 -53780
rect -160 -53940 -100 -53780
rect -380 -54040 -100 -53940
<< via3 >>
rect 900 2660 1100 2860
rect 1080 -25320 1360 -25120
<< metal4 >>
rect 800 3000 5400 3200
rect 800 2860 1200 3000
rect 800 2660 900 2860
rect 1100 2660 1200 2860
rect 800 2600 1200 2660
rect 1020 -25000 5340 -24800
rect 1020 -25120 1440 -25000
rect 1020 -25320 1080 -25120
rect 1360 -25320 1440 -25120
rect 1020 -25360 1440 -25320
use 2_to_4_decoder  2_to_4_decoder_0
timestamp 1671728743
transform 1 0 1060 0 1 -3080
box -460 -1920 2480 1848
use 3T  3T_0
timestamp 1671680485
transform 1 0 280 0 1 2300
box -280 -900 1153 838
use 3T  3T_1
timestamp 1671680485
transform 1 0 280 0 1 -53300
box -280 -900 1153 838
use 3T  3T_2
timestamp 1671680485
transform 1 0 480 0 1 -25700
box -280 -900 1153 838
use bias  bias_0
timestamp 1672278816
transform 1 0 17763 0 1 -60200
box 37 -200 5412 8450
use cd_current  cd_current_0
timestamp 1672331172
transform 1 0 1560 0 1 -54000
box 40 -200 5412 1200
use opamp_realcomp3_usefinger  opamp_realcomp3_usefinger_0
timestamp 1662739988
transform 1 0 5580 0 1 -60994
box -5380 594 6776 6403
use rc_model_4cap  rc_model_4cap_0
timestamp 1672330275
transform 1 0 -8000 0 1 19400
box 8000 -16400 25896 9200
use rc_model_6cap  rc_model_6cap_0
timestamp 1672329859
transform 1 0 -1400 0 1 -8600
box 1400 -16400 25896 9200
use rc_model_8cap  rc_model_8cap_0
timestamp 1672329920
transform 1 0 -1406 0 1 -36198
box 1400 -16400 25896 9200
use sample_hold  sample_hold_0
timestamp 1672262444
transform 1 0 7400 0 1 -60200
box 5200 -200 10099 4000
use sky130_fd_pr__pfet_01v8_lvt_BKTZ46  sky130_fd_pr__pfet_01v8_lvt_BKTZ46_0
timestamp 1672337038
transform 1 0 14757 0 1 -54334
box -957 -1866 957 1866
<< labels >>
flabel metal4 800 2860 1200 3200 0 FreeSans 1600 0 0 0 Vin_1
<< end >>
