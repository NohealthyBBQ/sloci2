magic
tech sky130A
magscale 1 2
timestamp 1672337919
<< metal1 >>
rect -960 3080 60 3100
rect -960 2980 -940 3080
rect -840 2980 60 3080
rect -960 2960 60 2980
rect 890 2660 900 2860
rect 1100 2660 1110 2860
rect -300 1700 300 1900
rect -960 -24920 360 -24900
rect -960 -25020 -940 -24920
rect -840 -25020 360 -24920
rect -960 -25040 360 -25020
rect -960 -52520 220 -52500
rect -960 -52620 -940 -52520
rect -840 -52620 220 -52520
rect -960 -52640 220 -52620
<< via1 >>
rect -940 2980 -840 3080
rect 900 2660 1100 2860
rect -940 -25020 -840 -24920
rect -940 -52620 -840 -52520
<< metal2 >>
rect -1000 3080 -800 3200
rect -1000 2980 -940 3080
rect -840 2980 -800 3080
rect -1000 -24920 -800 2980
rect 900 2860 1100 2870
rect 900 2650 1100 2660
rect -1000 -25020 -940 -24920
rect -840 -25020 -800 -24920
rect -1000 -52520 -800 -25020
rect -1000 -52620 -940 -52520
rect -840 -52620 -800 -52520
rect -1000 -52700 -800 -52620
<< via2 >>
rect 900 2660 1100 2860
<< metal3 >>
rect 890 2860 1110 2865
rect 890 2660 900 2860
rect 1100 2660 1110 2860
rect 890 2655 1110 2660
<< via3 >>
rect 900 2660 1100 2860
<< metal4 >>
rect 800 3000 5400 3200
rect 800 2860 1200 3000
rect 800 2660 900 2860
rect 1100 2660 1200 2860
rect 800 2600 1200 2660
use 2_to_4_decoder  2_to_4_decoder_0
timestamp 1671728743
transform 1 0 1060 0 1 -3080
box -460 -1920 2480 1848
use 3T  3T_0
timestamp 1671680485
transform 1 0 280 0 1 2300
box -280 -900 1153 838
use 3T  3T_1
timestamp 1671680485
transform 1 0 280 0 1 -53300
box -280 -900 1153 838
use 3T  3T_2
timestamp 1671680485
transform 1 0 480 0 1 -25700
box -280 -900 1153 838
use bias  bias_0
timestamp 1672278816
transform 1 0 17763 0 1 -60200
box 37 -200 5412 8450
use cd_current  cd_current_0
timestamp 1672331172
transform 1 0 1560 0 1 -54000
box 40 -200 5412 1200
use opamp_realcomp3_usefinger  opamp_realcomp3_usefinger_0
timestamp 1662739988
transform 1 0 5580 0 1 -60994
box -5380 594 6776 6403
use rc_model_4cap  rc_model_4cap_0
timestamp 1672330275
transform 1 0 -8000 0 1 19400
box 8000 -16400 25896 9200
use rc_model_6cap  rc_model_6cap_0
timestamp 1672329859
transform 1 0 -1400 0 1 -8600
box 1400 -16400 25896 9200
use rc_model_8cap  rc_model_8cap_0
timestamp 1672329920
transform 1 0 -1406 0 1 -36198
box 1400 -16400 25896 9200
use sample_hold  sample_hold_0
timestamp 1672262444
transform 1 0 7400 0 1 -60200
box 5200 -200 10099 4000
use sky130_fd_pr__pfet_01v8_lvt_BKTZ46  sky130_fd_pr__pfet_01v8_lvt_BKTZ46_0
timestamp 1672337038
transform 1 0 14757 0 1 -54334
box -957 -1866 957 1866
<< end >>
