magic
tech sky130A
magscale 1 2
timestamp 1662478139
<< pwell >>
rect -396 -519 396 519
<< nmoslvt >>
rect -200 109 200 309
rect -200 -309 200 -109
<< ndiff >>
rect -258 297 -200 309
rect -258 121 -246 297
rect -212 121 -200 297
rect -258 109 -200 121
rect 200 297 258 309
rect 200 121 212 297
rect 246 121 258 297
rect 200 109 258 121
rect -258 -121 -200 -109
rect -258 -297 -246 -121
rect -212 -297 -200 -121
rect -258 -309 -200 -297
rect 200 -121 258 -109
rect 200 -297 212 -121
rect 246 -297 258 -121
rect 200 -309 258 -297
<< ndiffc >>
rect -246 121 -212 297
rect 212 121 246 297
rect -246 -297 -212 -121
rect 212 -297 246 -121
<< psubdiff >>
rect -360 449 -264 483
rect 264 449 360 483
rect -360 387 -326 449
rect 326 387 360 449
rect -360 -449 -326 -387
rect 326 -449 360 -387
rect -360 -483 -264 -449
rect 264 -483 360 -449
<< psubdiffcont >>
rect -264 449 264 483
rect -360 -387 -326 387
rect 326 -387 360 387
rect -264 -483 264 -449
<< poly >>
rect -200 381 200 397
rect -200 347 -184 381
rect 184 347 200 381
rect -200 309 200 347
rect -200 71 200 109
rect -200 37 -184 71
rect 184 37 200 71
rect -200 21 200 37
rect -200 -37 200 -21
rect -200 -71 -184 -37
rect 184 -71 200 -37
rect -200 -109 200 -71
rect -200 -347 200 -309
rect -200 -381 -184 -347
rect 184 -381 200 -347
rect -200 -397 200 -381
<< polycont >>
rect -184 347 184 381
rect -184 37 184 71
rect -184 -71 184 -37
rect -184 -381 184 -347
<< locali >>
rect -360 449 -264 483
rect 264 449 360 483
rect -360 387 -326 449
rect 326 387 360 449
rect -200 347 -184 381
rect 184 347 200 381
rect -246 297 -212 313
rect -246 105 -212 121
rect 212 297 246 313
rect 212 105 246 121
rect -200 37 -184 71
rect 184 37 200 71
rect -200 -71 -184 -37
rect 184 -71 200 -37
rect -246 -121 -212 -105
rect -246 -313 -212 -297
rect 212 -121 246 -105
rect 212 -313 246 -297
rect -200 -381 -184 -347
rect 184 -381 200 -347
rect -360 -449 -326 -387
rect 326 -449 360 -387
rect -360 -483 -264 -449
rect 264 -483 360 -449
<< viali >>
rect -184 347 184 381
rect -246 121 -212 297
rect 212 121 246 297
rect -184 37 184 71
rect -184 -71 184 -37
rect -246 -297 -212 -121
rect 212 -297 246 -121
rect -184 -381 184 -347
<< metal1 >>
rect -196 381 196 387
rect -196 347 -184 381
rect 184 347 196 381
rect -196 341 196 347
rect -252 297 -206 309
rect -252 121 -246 297
rect -212 121 -206 297
rect -252 109 -206 121
rect 206 297 252 309
rect 206 121 212 297
rect 246 121 252 297
rect 206 109 252 121
rect -196 71 196 77
rect -196 37 -184 71
rect 184 37 196 71
rect -196 31 196 37
rect -196 -37 196 -31
rect -196 -71 -184 -37
rect 184 -71 196 -37
rect -196 -77 196 -71
rect -252 -121 -206 -109
rect -252 -297 -246 -121
rect -212 -297 -206 -121
rect -252 -309 -206 -297
rect 206 -121 252 -109
rect 206 -297 212 -121
rect 246 -297 252 -121
rect 206 -309 252 -297
rect -196 -347 196 -341
rect -196 -381 -184 -347
rect 184 -381 196 -347
rect -196 -387 196 -381
<< properties >>
string FIXED_BBOX -343 -466 343 466
string gencell sky130_fd_pr__nfet_01v8_lvt
string library sky130
string parameters w 1.0 l 2.0 m 2 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
