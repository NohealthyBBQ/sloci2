magic
tech sky130A
timestamp 1671827388
<< pwell >>
rect -564 -155 563 155
<< nmoslvt >>
rect -464 -50 -449 50
rect -416 -50 -401 50
rect -368 -50 -353 50
rect -320 -50 -305 50
rect -272 -50 -257 50
rect -224 -50 -209 50
rect -176 -50 -161 50
rect -128 -50 -113 50
rect -80 -50 -65 50
rect -32 -50 -17 50
rect 16 -50 31 50
rect 64 -50 79 50
rect 112 -50 127 50
rect 160 -50 175 50
rect 208 -50 223 50
rect 256 -50 271 50
rect 304 -50 319 50
rect 352 -50 367 50
rect 400 -50 415 50
rect 448 -50 463 50
<< ndiff >>
rect -495 44 -464 50
rect -495 -44 -489 44
rect -472 -44 -464 44
rect -495 -50 -464 -44
rect -449 44 -416 50
rect -449 -44 -441 44
rect -424 -44 -416 44
rect -449 -50 -416 -44
rect -401 44 -368 50
rect -401 -44 -393 44
rect -376 -44 -368 44
rect -401 -50 -368 -44
rect -353 44 -320 50
rect -353 -44 -345 44
rect -328 -44 -320 44
rect -353 -50 -320 -44
rect -305 44 -272 50
rect -305 -44 -297 44
rect -280 -44 -272 44
rect -305 -50 -272 -44
rect -257 44 -224 50
rect -257 -44 -249 44
rect -232 -44 -224 44
rect -257 -50 -224 -44
rect -209 44 -176 50
rect -209 -44 -201 44
rect -184 -44 -176 44
rect -209 -50 -176 -44
rect -161 44 -128 50
rect -161 -44 -153 44
rect -136 -44 -128 44
rect -161 -50 -128 -44
rect -113 44 -80 50
rect -113 -44 -105 44
rect -88 -44 -80 44
rect -113 -50 -80 -44
rect -65 44 -32 50
rect -65 -44 -57 44
rect -40 -44 -32 44
rect -65 -50 -32 -44
rect -17 44 16 50
rect -17 -44 -9 44
rect 8 -44 16 44
rect -17 -50 16 -44
rect 31 44 64 50
rect 31 -44 39 44
rect 56 -44 64 44
rect 31 -50 64 -44
rect 79 44 112 50
rect 79 -44 87 44
rect 104 -44 112 44
rect 79 -50 112 -44
rect 127 44 160 50
rect 127 -44 135 44
rect 152 -44 160 44
rect 127 -50 160 -44
rect 175 44 208 50
rect 175 -44 183 44
rect 200 -44 208 44
rect 175 -50 208 -44
rect 223 44 256 50
rect 223 -44 231 44
rect 248 -44 256 44
rect 223 -50 256 -44
rect 271 44 304 50
rect 271 -44 279 44
rect 296 -44 304 44
rect 271 -50 304 -44
rect 319 44 352 50
rect 319 -44 327 44
rect 344 -44 352 44
rect 319 -50 352 -44
rect 367 44 400 50
rect 367 -44 375 44
rect 392 -44 400 44
rect 367 -50 400 -44
rect 415 44 448 50
rect 415 -44 423 44
rect 440 -44 448 44
rect 415 -50 448 -44
rect 463 44 494 50
rect 463 -44 471 44
rect 488 -44 494 44
rect 463 -50 494 -44
<< ndiffc >>
rect -489 -44 -472 44
rect -441 -44 -424 44
rect -393 -44 -376 44
rect -345 -44 -328 44
rect -297 -44 -280 44
rect -249 -44 -232 44
rect -201 -44 -184 44
rect -153 -44 -136 44
rect -105 -44 -88 44
rect -57 -44 -40 44
rect -9 -44 8 44
rect 39 -44 56 44
rect 87 -44 104 44
rect 135 -44 152 44
rect 183 -44 200 44
rect 231 -44 248 44
rect 279 -44 296 44
rect 327 -44 344 44
rect 375 -44 392 44
rect 423 -44 440 44
rect 471 -44 488 44
<< psubdiff >>
rect -546 120 -498 137
rect 497 120 545 137
rect -546 89 -529 120
rect 528 89 545 120
rect -546 -120 -529 -89
rect 528 -120 545 -89
rect -546 -137 -498 -120
rect 497 -137 545 -120
<< psubdiffcont >>
rect -498 120 497 137
rect -546 -89 -529 89
rect 528 -89 545 89
rect -498 -137 497 -120
<< poly >>
rect -464 50 -449 63
rect -416 50 -401 63
rect -368 50 -353 63
rect -320 50 -305 63
rect -272 50 -257 63
rect -224 50 -209 63
rect -176 50 -161 63
rect -128 50 -113 63
rect -80 50 -65 63
rect -32 50 -17 63
rect 16 50 31 63
rect 64 50 79 63
rect 112 50 127 63
rect 160 50 175 63
rect 208 50 223 63
rect 256 50 271 63
rect 304 50 319 63
rect 352 50 367 63
rect 400 50 415 63
rect 448 50 463 63
rect -464 -61 -449 -50
rect -416 -61 -401 -50
rect -368 -61 -353 -50
rect -320 -61 -305 -50
rect -272 -61 -257 -50
rect -224 -61 -209 -50
rect -176 -61 -161 -50
rect -128 -61 -113 -50
rect -80 -61 -65 -50
rect -32 -61 -17 -50
rect 16 -61 31 -50
rect 64 -61 79 -50
rect 112 -61 127 -50
rect 160 -61 175 -50
rect 208 -61 223 -50
rect 256 -61 271 -50
rect 304 -61 319 -50
rect 352 -61 367 -50
rect 400 -61 415 -50
rect 448 -61 463 -50
rect -473 -69 463 -61
rect -473 -86 15 -69
rect 32 -86 463 -69
rect -473 -94 -440 -86
rect -377 -94 -344 -86
rect -281 -94 -248 -86
rect -185 -94 -152 -86
rect -89 -94 -56 -86
rect 7 -94 40 -86
rect 103 -94 136 -86
rect 199 -94 232 -86
rect 295 -94 328 -86
rect 391 -94 424 -86
<< polycont >>
rect 15 -86 32 -69
<< locali >>
rect -546 120 -498 137
rect 497 120 545 137
rect -546 89 -529 120
rect 528 89 545 120
rect -489 44 -472 52
rect -489 -52 -472 -44
rect -441 44 -424 52
rect -441 -52 -424 -44
rect -393 44 -376 52
rect -393 -52 -376 -44
rect -345 44 -328 52
rect -345 -52 -328 -44
rect -297 44 -280 52
rect -297 -52 -280 -44
rect -249 44 -232 52
rect -249 -52 -232 -44
rect -201 44 -184 52
rect -201 -52 -184 -44
rect -153 44 -136 52
rect -153 -52 -136 -44
rect -105 44 -88 52
rect -105 -52 -88 -44
rect -57 44 -40 52
rect -57 -52 -40 -44
rect -9 44 8 52
rect -9 -52 8 -44
rect 39 44 56 52
rect 39 -52 56 -44
rect 87 44 104 52
rect 87 -52 104 -44
rect 135 44 152 52
rect 135 -52 152 -44
rect 183 44 200 52
rect 183 -52 200 -44
rect 231 44 248 52
rect 231 -52 248 -44
rect 279 44 296 52
rect 279 -52 296 -44
rect 327 44 344 52
rect 327 -52 344 -44
rect 375 44 392 52
rect 375 -52 392 -44
rect 423 44 440 52
rect 423 -52 440 -44
rect 471 44 488 52
rect 471 -52 488 -44
rect 7 -86 15 -69
rect 32 -86 40 -69
rect -546 -120 -529 -89
rect 528 -120 545 -89
rect -546 -137 -498 -120
rect 497 -137 545 -120
<< viali >>
rect -489 -44 -472 44
rect -441 -44 -424 44
rect -393 -44 -376 44
rect -345 -44 -328 44
rect -297 -44 -280 44
rect -249 -44 -232 44
rect -201 -44 -184 44
rect -153 -44 -136 44
rect -105 -44 -88 44
rect -57 -44 -40 44
rect -9 -44 8 44
rect 39 -44 56 44
rect 87 -44 104 44
rect 135 -44 152 44
rect 183 -44 200 44
rect 231 -44 248 44
rect 279 -44 296 44
rect 327 -44 344 44
rect 375 -44 392 44
rect 423 -44 440 44
rect 471 -44 488 44
rect 15 -86 32 -69
<< metal1 >>
rect -492 44 -469 50
rect -492 -14 -489 44
rect -497 -17 -489 -14
rect -472 -14 -469 44
rect -449 47 -416 50
rect -449 17 -445 47
rect -419 17 -416 47
rect -449 14 -441 17
rect -472 -17 -464 -14
rect -497 -47 -493 -17
rect -467 -47 -464 -17
rect -497 -50 -464 -47
rect -444 -44 -441 14
rect -424 14 -416 17
rect -396 44 -373 50
rect -424 -44 -421 14
rect -396 -14 -393 44
rect -444 -50 -421 -44
rect -401 -17 -393 -14
rect -376 -14 -373 44
rect -353 47 -320 50
rect -353 17 -349 47
rect -323 17 -320 47
rect -353 14 -345 17
rect -376 -17 -368 -14
rect -401 -47 -397 -17
rect -371 -47 -368 -17
rect -401 -50 -368 -47
rect -348 -44 -345 14
rect -328 14 -320 17
rect -300 44 -277 50
rect -328 -44 -325 14
rect -300 -14 -297 44
rect -348 -50 -325 -44
rect -305 -17 -297 -14
rect -280 -14 -277 44
rect -257 47 -224 50
rect -257 17 -253 47
rect -227 17 -224 47
rect -257 14 -249 17
rect -280 -17 -272 -14
rect -305 -47 -301 -17
rect -275 -47 -272 -17
rect -305 -50 -272 -47
rect -252 -44 -249 14
rect -232 14 -224 17
rect -204 44 -181 50
rect -232 -44 -229 14
rect -204 -14 -201 44
rect -252 -50 -229 -44
rect -209 -17 -201 -14
rect -184 -14 -181 44
rect -161 47 -128 50
rect -161 17 -157 47
rect -131 17 -128 47
rect -161 14 -153 17
rect -184 -17 -176 -14
rect -209 -47 -205 -17
rect -179 -47 -176 -17
rect -209 -50 -176 -47
rect -156 -44 -153 14
rect -136 14 -128 17
rect -108 44 -85 50
rect -136 -44 -133 14
rect -108 -14 -105 44
rect -156 -50 -133 -44
rect -113 -17 -105 -14
rect -88 -14 -85 44
rect -65 47 -32 50
rect -65 17 -61 47
rect -35 17 -32 47
rect -65 14 -57 17
rect -88 -17 -80 -14
rect -113 -47 -109 -17
rect -83 -47 -80 -17
rect -113 -50 -80 -47
rect -60 -44 -57 14
rect -40 14 -32 17
rect -12 44 11 50
rect -40 -44 -37 14
rect -12 -14 -9 44
rect -60 -50 -37 -44
rect -17 -17 -9 -14
rect 8 -14 11 44
rect 31 47 64 50
rect 31 17 35 47
rect 61 17 64 47
rect 31 14 39 17
rect 8 -17 16 -14
rect -17 -47 -13 -17
rect 13 -47 16 -17
rect -17 -50 16 -47
rect 36 -44 39 14
rect 56 14 64 17
rect 84 44 107 50
rect 56 -44 59 14
rect 84 -14 87 44
rect 36 -50 59 -44
rect 79 -17 87 -14
rect 104 -14 107 44
rect 127 47 160 50
rect 127 17 131 47
rect 157 17 160 47
rect 127 14 135 17
rect 104 -17 112 -14
rect 79 -47 83 -17
rect 109 -47 112 -17
rect 79 -50 112 -47
rect 132 -44 135 14
rect 152 14 160 17
rect 180 44 203 50
rect 152 -44 155 14
rect 180 -14 183 44
rect 132 -50 155 -44
rect 175 -17 183 -14
rect 200 -14 203 44
rect 223 47 256 50
rect 223 17 227 47
rect 253 17 256 47
rect 223 14 231 17
rect 200 -17 208 -14
rect 175 -47 179 -17
rect 205 -47 208 -17
rect 175 -50 208 -47
rect 228 -44 231 14
rect 248 14 256 17
rect 276 44 299 50
rect 248 -44 251 14
rect 276 -14 279 44
rect 228 -50 251 -44
rect 271 -17 279 -14
rect 296 -14 299 44
rect 319 47 352 50
rect 319 17 323 47
rect 349 17 352 47
rect 319 14 327 17
rect 296 -17 304 -14
rect 271 -47 275 -17
rect 301 -47 304 -17
rect 271 -50 304 -47
rect 324 -44 327 14
rect 344 14 352 17
rect 372 44 395 50
rect 344 -44 347 14
rect 372 -14 375 44
rect 324 -50 347 -44
rect 367 -17 375 -14
rect 392 -14 395 44
rect 415 47 448 50
rect 415 17 419 47
rect 445 17 448 47
rect 415 14 423 17
rect 392 -17 400 -14
rect 367 -47 371 -17
rect 397 -47 400 -17
rect 367 -50 400 -47
rect 420 -44 423 14
rect 440 14 448 17
rect 468 44 491 50
rect 440 -44 443 14
rect 468 -14 471 44
rect 420 -50 443 -44
rect 463 -17 471 -14
rect 488 -14 491 44
rect 488 -17 496 -14
rect 463 -47 467 -17
rect 493 -47 496 -17
rect 463 -50 496 -47
rect -473 -69 463 -66
rect -473 -86 15 -69
rect 32 -86 463 -69
rect -473 -90 463 -86
<< via1 >>
rect -445 44 -419 47
rect -445 17 -441 44
rect -441 17 -424 44
rect -424 17 -419 44
rect -493 -44 -489 -17
rect -489 -44 -472 -17
rect -472 -44 -467 -17
rect -493 -47 -467 -44
rect -349 44 -323 47
rect -349 17 -345 44
rect -345 17 -328 44
rect -328 17 -323 44
rect -397 -44 -393 -17
rect -393 -44 -376 -17
rect -376 -44 -371 -17
rect -397 -47 -371 -44
rect -253 44 -227 47
rect -253 17 -249 44
rect -249 17 -232 44
rect -232 17 -227 44
rect -301 -44 -297 -17
rect -297 -44 -280 -17
rect -280 -44 -275 -17
rect -301 -47 -275 -44
rect -157 44 -131 47
rect -157 17 -153 44
rect -153 17 -136 44
rect -136 17 -131 44
rect -205 -44 -201 -17
rect -201 -44 -184 -17
rect -184 -44 -179 -17
rect -205 -47 -179 -44
rect -61 44 -35 47
rect -61 17 -57 44
rect -57 17 -40 44
rect -40 17 -35 44
rect -109 -44 -105 -17
rect -105 -44 -88 -17
rect -88 -44 -83 -17
rect -109 -47 -83 -44
rect 35 44 61 47
rect 35 17 39 44
rect 39 17 56 44
rect 56 17 61 44
rect -13 -44 -9 -17
rect -9 -44 8 -17
rect 8 -44 13 -17
rect -13 -47 13 -44
rect 131 44 157 47
rect 131 17 135 44
rect 135 17 152 44
rect 152 17 157 44
rect 83 -44 87 -17
rect 87 -44 104 -17
rect 104 -44 109 -17
rect 83 -47 109 -44
rect 227 44 253 47
rect 227 17 231 44
rect 231 17 248 44
rect 248 17 253 44
rect 179 -44 183 -17
rect 183 -44 200 -17
rect 200 -44 205 -17
rect 179 -47 205 -44
rect 323 44 349 47
rect 323 17 327 44
rect 327 17 344 44
rect 344 17 349 44
rect 275 -44 279 -17
rect 279 -44 296 -17
rect 296 -44 301 -17
rect 275 -47 301 -44
rect 419 44 445 47
rect 419 17 423 44
rect 423 17 440 44
rect 440 17 445 44
rect 371 -44 375 -17
rect 375 -44 392 -17
rect 392 -44 397 -17
rect 371 -47 397 -44
rect 467 -44 471 -17
rect 471 -44 488 -17
rect 488 -44 493 -17
rect 467 -47 493 -44
<< metal2 >>
rect -497 47 498 94
rect -497 17 -445 47
rect -419 17 -349 47
rect -323 17 -253 47
rect -227 17 -157 47
rect -131 17 -61 47
rect -35 17 35 47
rect 61 17 131 47
rect 157 17 227 47
rect 253 17 323 47
rect 349 17 419 47
rect 445 17 498 47
rect -497 14 498 17
rect -498 -17 497 -14
rect -498 -47 -493 -17
rect -467 -47 -397 -17
rect -371 -47 -301 -17
rect -275 -47 -205 -17
rect -179 -47 -109 -17
rect -83 -47 -13 -17
rect 13 -47 83 -17
rect 109 -47 179 -17
rect 205 -47 275 -17
rect 301 -47 371 -17
rect 397 -47 467 -17
rect 493 -47 497 -17
rect -498 -94 497 -47
<< properties >>
string FIXED_BBOX -537 -128 537 128
string gencell sky130_fd_pr__nfet_01v8_lvt
string library sky130
string parameters w 1.0 l 0.15 m 1 nf 20 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
