magic
tech sky130A
magscale 1 2
timestamp 1662404926
<< error_p >>
rect -607 181 -545 187
rect -479 181 -417 187
rect -351 181 -289 187
rect -223 181 -161 187
rect -95 181 -33 187
rect 33 181 95 187
rect 161 181 223 187
rect 289 181 351 187
rect 417 181 479 187
rect 545 181 607 187
rect -607 147 -595 181
rect -479 147 -467 181
rect -351 147 -339 181
rect -223 147 -211 181
rect -95 147 -83 181
rect 33 147 45 181
rect 161 147 173 181
rect 289 147 301 181
rect 417 147 429 181
rect 545 147 557 181
rect -607 141 -545 147
rect -479 141 -417 147
rect -351 141 -289 147
rect -223 141 -161 147
rect -95 141 -33 147
rect 33 141 95 147
rect 161 141 223 147
rect 289 141 351 147
rect 417 141 479 147
rect 545 141 607 147
rect -607 -147 -545 -141
rect -479 -147 -417 -141
rect -351 -147 -289 -141
rect -223 -147 -161 -141
rect -95 -147 -33 -141
rect 33 -147 95 -141
rect 161 -147 223 -141
rect 289 -147 351 -141
rect 417 -147 479 -141
rect 545 -147 607 -141
rect -607 -181 -595 -147
rect -479 -181 -467 -147
rect -351 -181 -339 -147
rect -223 -181 -211 -147
rect -95 -181 -83 -147
rect 33 -181 45 -147
rect 161 -181 173 -147
rect 289 -181 301 -147
rect 417 -181 429 -147
rect 545 -181 557 -147
rect -607 -187 -545 -181
rect -479 -187 -417 -181
rect -351 -187 -289 -181
rect -223 -187 -161 -181
rect -95 -187 -33 -181
rect 33 -187 95 -181
rect 161 -187 223 -181
rect 289 -187 351 -181
rect 417 -187 479 -181
rect 545 -187 607 -181
<< nwell >>
rect -807 -319 807 319
<< pmoslvt >>
rect -611 -100 -541 100
rect -483 -100 -413 100
rect -355 -100 -285 100
rect -227 -100 -157 100
rect -99 -100 -29 100
rect 29 -100 99 100
rect 157 -100 227 100
rect 285 -100 355 100
rect 413 -100 483 100
rect 541 -100 611 100
<< pdiff >>
rect -669 88 -611 100
rect -669 -88 -657 88
rect -623 -88 -611 88
rect -669 -100 -611 -88
rect -541 88 -483 100
rect -541 -88 -529 88
rect -495 -88 -483 88
rect -541 -100 -483 -88
rect -413 88 -355 100
rect -413 -88 -401 88
rect -367 -88 -355 88
rect -413 -100 -355 -88
rect -285 88 -227 100
rect -285 -88 -273 88
rect -239 -88 -227 88
rect -285 -100 -227 -88
rect -157 88 -99 100
rect -157 -88 -145 88
rect -111 -88 -99 88
rect -157 -100 -99 -88
rect -29 88 29 100
rect -29 -88 -17 88
rect 17 -88 29 88
rect -29 -100 29 -88
rect 99 88 157 100
rect 99 -88 111 88
rect 145 -88 157 88
rect 99 -100 157 -88
rect 227 88 285 100
rect 227 -88 239 88
rect 273 -88 285 88
rect 227 -100 285 -88
rect 355 88 413 100
rect 355 -88 367 88
rect 401 -88 413 88
rect 355 -100 413 -88
rect 483 88 541 100
rect 483 -88 495 88
rect 529 -88 541 88
rect 483 -100 541 -88
rect 611 88 669 100
rect 611 -88 623 88
rect 657 -88 669 88
rect 611 -100 669 -88
<< pdiffc >>
rect -657 -88 -623 88
rect -529 -88 -495 88
rect -401 -88 -367 88
rect -273 -88 -239 88
rect -145 -88 -111 88
rect -17 -88 17 88
rect 111 -88 145 88
rect 239 -88 273 88
rect 367 -88 401 88
rect 495 -88 529 88
rect 623 -88 657 88
<< nsubdiff >>
rect -771 249 -675 283
rect 675 249 771 283
rect -771 187 -737 249
rect 737 187 771 249
rect -771 -249 -737 -187
rect 737 -249 771 -187
rect -771 -283 -675 -249
rect 675 -283 771 -249
<< nsubdiffcont >>
rect -675 249 675 283
rect -771 -187 -737 187
rect 737 -187 771 187
rect -675 -283 675 -249
<< poly >>
rect -611 181 -541 197
rect -611 147 -595 181
rect -557 147 -541 181
rect -611 100 -541 147
rect -483 181 -413 197
rect -483 147 -467 181
rect -429 147 -413 181
rect -483 100 -413 147
rect -355 181 -285 197
rect -355 147 -339 181
rect -301 147 -285 181
rect -355 100 -285 147
rect -227 181 -157 197
rect -227 147 -211 181
rect -173 147 -157 181
rect -227 100 -157 147
rect -99 181 -29 197
rect -99 147 -83 181
rect -45 147 -29 181
rect -99 100 -29 147
rect 29 181 99 197
rect 29 147 45 181
rect 83 147 99 181
rect 29 100 99 147
rect 157 181 227 197
rect 157 147 173 181
rect 211 147 227 181
rect 157 100 227 147
rect 285 181 355 197
rect 285 147 301 181
rect 339 147 355 181
rect 285 100 355 147
rect 413 181 483 197
rect 413 147 429 181
rect 467 147 483 181
rect 413 100 483 147
rect 541 181 611 197
rect 541 147 557 181
rect 595 147 611 181
rect 541 100 611 147
rect -611 -147 -541 -100
rect -611 -181 -595 -147
rect -557 -181 -541 -147
rect -611 -197 -541 -181
rect -483 -147 -413 -100
rect -483 -181 -467 -147
rect -429 -181 -413 -147
rect -483 -197 -413 -181
rect -355 -147 -285 -100
rect -355 -181 -339 -147
rect -301 -181 -285 -147
rect -355 -197 -285 -181
rect -227 -147 -157 -100
rect -227 -181 -211 -147
rect -173 -181 -157 -147
rect -227 -197 -157 -181
rect -99 -147 -29 -100
rect -99 -181 -83 -147
rect -45 -181 -29 -147
rect -99 -197 -29 -181
rect 29 -147 99 -100
rect 29 -181 45 -147
rect 83 -181 99 -147
rect 29 -197 99 -181
rect 157 -147 227 -100
rect 157 -181 173 -147
rect 211 -181 227 -147
rect 157 -197 227 -181
rect 285 -147 355 -100
rect 285 -181 301 -147
rect 339 -181 355 -147
rect 285 -197 355 -181
rect 413 -147 483 -100
rect 413 -181 429 -147
rect 467 -181 483 -147
rect 413 -197 483 -181
rect 541 -147 611 -100
rect 541 -181 557 -147
rect 595 -181 611 -147
rect 541 -197 611 -181
<< polycont >>
rect -595 147 -557 181
rect -467 147 -429 181
rect -339 147 -301 181
rect -211 147 -173 181
rect -83 147 -45 181
rect 45 147 83 181
rect 173 147 211 181
rect 301 147 339 181
rect 429 147 467 181
rect 557 147 595 181
rect -595 -181 -557 -147
rect -467 -181 -429 -147
rect -339 -181 -301 -147
rect -211 -181 -173 -147
rect -83 -181 -45 -147
rect 45 -181 83 -147
rect 173 -181 211 -147
rect 301 -181 339 -147
rect 429 -181 467 -147
rect 557 -181 595 -147
<< locali >>
rect -771 249 -675 283
rect 675 249 771 283
rect -771 187 -737 249
rect 737 187 771 249
rect -611 147 -595 181
rect -557 147 -541 181
rect -483 147 -467 181
rect -429 147 -413 181
rect -355 147 -339 181
rect -301 147 -285 181
rect -227 147 -211 181
rect -173 147 -157 181
rect -99 147 -83 181
rect -45 147 -29 181
rect 29 147 45 181
rect 83 147 99 181
rect 157 147 173 181
rect 211 147 227 181
rect 285 147 301 181
rect 339 147 355 181
rect 413 147 429 181
rect 467 147 483 181
rect 541 147 557 181
rect 595 147 611 181
rect -657 88 -623 104
rect -657 -104 -623 -88
rect -529 88 -495 104
rect -529 -104 -495 -88
rect -401 88 -367 104
rect -401 -104 -367 -88
rect -273 88 -239 104
rect -273 -104 -239 -88
rect -145 88 -111 104
rect -145 -104 -111 -88
rect -17 88 17 104
rect -17 -104 17 -88
rect 111 88 145 104
rect 111 -104 145 -88
rect 239 88 273 104
rect 239 -104 273 -88
rect 367 88 401 104
rect 367 -104 401 -88
rect 495 88 529 104
rect 495 -104 529 -88
rect 623 88 657 104
rect 623 -104 657 -88
rect -611 -181 -595 -147
rect -557 -181 -541 -147
rect -483 -181 -467 -147
rect -429 -181 -413 -147
rect -355 -181 -339 -147
rect -301 -181 -285 -147
rect -227 -181 -211 -147
rect -173 -181 -157 -147
rect -99 -181 -83 -147
rect -45 -181 -29 -147
rect 29 -181 45 -147
rect 83 -181 99 -147
rect 157 -181 173 -147
rect 211 -181 227 -147
rect 285 -181 301 -147
rect 339 -181 355 -147
rect 413 -181 429 -147
rect 467 -181 483 -147
rect 541 -181 557 -147
rect 595 -181 611 -147
rect -771 -249 -737 -187
rect 737 -249 771 -187
rect -771 -283 -675 -249
rect 675 -283 771 -249
<< viali >>
rect -595 147 -557 181
rect -467 147 -429 181
rect -339 147 -301 181
rect -211 147 -173 181
rect -83 147 -45 181
rect 45 147 83 181
rect 173 147 211 181
rect 301 147 339 181
rect 429 147 467 181
rect 557 147 595 181
rect -657 -88 -623 88
rect -529 -88 -495 88
rect -401 -88 -367 88
rect -273 -88 -239 88
rect -145 -88 -111 88
rect -17 -88 17 88
rect 111 -88 145 88
rect 239 -88 273 88
rect 367 -88 401 88
rect 495 -88 529 88
rect 623 -88 657 88
rect -595 -181 -557 -147
rect -467 -181 -429 -147
rect -339 -181 -301 -147
rect -211 -181 -173 -147
rect -83 -181 -45 -147
rect 45 -181 83 -147
rect 173 -181 211 -147
rect 301 -181 339 -147
rect 429 -181 467 -147
rect 557 -181 595 -147
<< metal1 >>
rect -607 181 -545 187
rect -607 147 -595 181
rect -557 147 -545 181
rect -607 141 -545 147
rect -479 181 -417 187
rect -479 147 -467 181
rect -429 147 -417 181
rect -479 141 -417 147
rect -351 181 -289 187
rect -351 147 -339 181
rect -301 147 -289 181
rect -351 141 -289 147
rect -223 181 -161 187
rect -223 147 -211 181
rect -173 147 -161 181
rect -223 141 -161 147
rect -95 181 -33 187
rect -95 147 -83 181
rect -45 147 -33 181
rect -95 141 -33 147
rect 33 181 95 187
rect 33 147 45 181
rect 83 147 95 181
rect 33 141 95 147
rect 161 181 223 187
rect 161 147 173 181
rect 211 147 223 181
rect 161 141 223 147
rect 289 181 351 187
rect 289 147 301 181
rect 339 147 351 181
rect 289 141 351 147
rect 417 181 479 187
rect 417 147 429 181
rect 467 147 479 181
rect 417 141 479 147
rect 545 181 607 187
rect 545 147 557 181
rect 595 147 607 181
rect 545 141 607 147
rect -663 88 -617 100
rect -663 -88 -657 88
rect -623 -88 -617 88
rect -663 -100 -617 -88
rect -535 88 -489 100
rect -535 -88 -529 88
rect -495 -88 -489 88
rect -535 -100 -489 -88
rect -407 88 -361 100
rect -407 -88 -401 88
rect -367 -88 -361 88
rect -407 -100 -361 -88
rect -279 88 -233 100
rect -279 -88 -273 88
rect -239 -88 -233 88
rect -279 -100 -233 -88
rect -151 88 -105 100
rect -151 -88 -145 88
rect -111 -88 -105 88
rect -151 -100 -105 -88
rect -23 88 23 100
rect -23 -88 -17 88
rect 17 -88 23 88
rect -23 -100 23 -88
rect 105 88 151 100
rect 105 -88 111 88
rect 145 -88 151 88
rect 105 -100 151 -88
rect 233 88 279 100
rect 233 -88 239 88
rect 273 -88 279 88
rect 233 -100 279 -88
rect 361 88 407 100
rect 361 -88 367 88
rect 401 -88 407 88
rect 361 -100 407 -88
rect 489 88 535 100
rect 489 -88 495 88
rect 529 -88 535 88
rect 489 -100 535 -88
rect 617 88 663 100
rect 617 -88 623 88
rect 657 -88 663 88
rect 617 -100 663 -88
rect -607 -147 -545 -141
rect -607 -181 -595 -147
rect -557 -181 -545 -147
rect -607 -187 -545 -181
rect -479 -147 -417 -141
rect -479 -181 -467 -147
rect -429 -181 -417 -147
rect -479 -187 -417 -181
rect -351 -147 -289 -141
rect -351 -181 -339 -147
rect -301 -181 -289 -147
rect -351 -187 -289 -181
rect -223 -147 -161 -141
rect -223 -181 -211 -147
rect -173 -181 -161 -147
rect -223 -187 -161 -181
rect -95 -147 -33 -141
rect -95 -181 -83 -147
rect -45 -181 -33 -147
rect -95 -187 -33 -181
rect 33 -147 95 -141
rect 33 -181 45 -147
rect 83 -181 95 -147
rect 33 -187 95 -181
rect 161 -147 223 -141
rect 161 -181 173 -147
rect 211 -181 223 -147
rect 161 -187 223 -181
rect 289 -147 351 -141
rect 289 -181 301 -147
rect 339 -181 351 -147
rect 289 -187 351 -181
rect 417 -147 479 -141
rect 417 -181 429 -147
rect 467 -181 479 -147
rect 417 -187 479 -181
rect 545 -147 607 -141
rect 545 -181 557 -147
rect 595 -181 607 -147
rect 545 -187 607 -181
<< properties >>
string FIXED_BBOX -754 -266 754 266
string gencell sky130_fd_pr__pfet_01v8_lvt
string library sky130
string parameters w 1.0 l 0.35 m 1 nf 10 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.35 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
