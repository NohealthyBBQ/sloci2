magic
tech sky130A
magscale 1 2
timestamp 1662983156
<< error_p >>
rect -29 309 29 315
rect -29 275 -17 309
rect -29 269 29 275
rect -29 71 29 77
rect -29 37 -17 71
rect -29 31 29 37
rect -29 -37 29 -31
rect -29 -71 -17 -37
rect -29 -77 29 -71
rect -29 -275 29 -269
rect -29 -309 -17 -275
rect -29 -315 29 -309
<< pwell >>
rect -211 -447 211 447
<< nmoslvt >>
rect -15 109 15 237
rect -15 -237 15 -109
<< ndiff >>
rect -73 225 -15 237
rect -73 121 -61 225
rect -27 121 -15 225
rect -73 109 -15 121
rect 15 225 73 237
rect 15 121 27 225
rect 61 121 73 225
rect 15 109 73 121
rect -73 -121 -15 -109
rect -73 -225 -61 -121
rect -27 -225 -15 -121
rect -73 -237 -15 -225
rect 15 -121 73 -109
rect 15 -225 27 -121
rect 61 -225 73 -121
rect 15 -237 73 -225
<< ndiffc >>
rect -61 121 -27 225
rect 27 121 61 225
rect -61 -225 -27 -121
rect 27 -225 61 -121
<< psubdiff >>
rect -175 377 -79 411
rect 79 377 175 411
rect -175 315 -141 377
rect 141 315 175 377
rect -175 -377 -141 -315
rect 141 -377 175 -315
rect -175 -411 -79 -377
rect 79 -411 175 -377
<< psubdiffcont >>
rect -79 377 79 411
rect -175 -315 -141 315
rect 141 -315 175 315
rect -79 -411 79 -377
<< poly >>
rect -33 309 33 325
rect -33 275 -17 309
rect 17 275 33 309
rect -33 259 33 275
rect -15 237 15 259
rect -15 87 15 109
rect -33 71 33 87
rect -33 37 -17 71
rect 17 37 33 71
rect -33 21 33 37
rect -33 -37 33 -21
rect -33 -71 -17 -37
rect 17 -71 33 -37
rect -33 -87 33 -71
rect -15 -109 15 -87
rect -15 -259 15 -237
rect -33 -275 33 -259
rect -33 -309 -17 -275
rect 17 -309 33 -275
rect -33 -325 33 -309
<< polycont >>
rect -17 275 17 309
rect -17 37 17 71
rect -17 -71 17 -37
rect -17 -309 17 -275
<< locali >>
rect -175 377 -79 411
rect 79 377 175 411
rect -175 315 -141 377
rect 141 315 175 377
rect -33 275 -17 309
rect 17 275 33 309
rect -61 225 -27 241
rect -61 105 -27 121
rect 27 225 61 241
rect 27 105 61 121
rect -33 37 -17 71
rect 17 37 33 71
rect -33 -71 -17 -37
rect 17 -71 33 -37
rect -61 -121 -27 -105
rect -61 -241 -27 -225
rect 27 -121 61 -105
rect 27 -241 61 -225
rect -33 -309 -17 -275
rect 17 -309 33 -275
rect -175 -377 -141 -315
rect 141 -377 175 -315
rect -175 -411 -79 -377
rect 79 -411 175 -377
<< viali >>
rect -17 275 17 309
rect -61 121 -27 225
rect 27 121 61 225
rect -17 37 17 71
rect -17 -71 17 -37
rect -61 -225 -27 -121
rect 27 -225 61 -121
rect -17 -309 17 -275
<< metal1 >>
rect -29 309 29 315
rect -29 275 -17 309
rect 17 275 29 309
rect -29 269 29 275
rect -67 225 -21 237
rect -67 121 -61 225
rect -27 121 -21 225
rect -67 109 -21 121
rect 21 225 67 237
rect 21 121 27 225
rect 61 121 67 225
rect 21 109 67 121
rect -29 71 29 77
rect -29 37 -17 71
rect 17 37 29 71
rect -29 31 29 37
rect -29 -37 29 -31
rect -29 -71 -17 -37
rect 17 -71 29 -37
rect -29 -77 29 -71
rect -67 -121 -21 -109
rect -67 -225 -61 -121
rect -27 -225 -21 -121
rect -67 -237 -21 -225
rect 21 -121 67 -109
rect 21 -225 27 -121
rect 61 -225 67 -121
rect 21 -237 67 -225
rect -29 -275 29 -269
rect -29 -309 -17 -275
rect 17 -309 29 -275
rect -29 -315 29 -309
<< properties >>
string FIXED_BBOX -158 -394 158 394
string gencell sky130_fd_pr__nfet_01v8_lvt
string library sky130
string parameters w 0.64 l 0.150 m 2 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
