magic
tech sky130A
magscale 1 2
timestamp 1672331172
<< locali >>
rect 180 360 240 540
rect 1100 360 1160 540
rect 2020 360 2080 540
rect 2920 360 2980 540
rect 3840 360 3900 540
rect 4760 360 4820 540
rect 5220 360 5280 540
<< metal1 >>
rect 180 160 280 900
rect 1080 870 4380 900
rect 1070 700 1080 780
rect 1160 700 1170 780
rect 1990 700 2000 780
rect 2080 700 2090 780
rect 2910 700 2920 780
rect 3000 700 3010 780
rect 3810 700 3820 780
rect 3900 700 3910 780
rect 4730 700 4740 780
rect 4820 700 4830 780
rect 640 580 700 680
rect 1560 580 1620 680
rect 2480 580 2540 680
rect 3380 580 3440 680
rect 4300 580 4360 680
rect 640 480 4360 580
rect 640 380 700 480
rect 1560 380 1620 480
rect 2480 380 2540 480
rect 3380 380 3440 480
rect 4300 380 4360 480
rect 1080 160 4380 190
rect 5160 160 5280 920
<< via1 >>
rect 1080 700 1160 780
rect 2000 700 2080 780
rect 2920 700 3000 780
rect 3820 700 3900 780
rect 4740 700 4820 780
<< metal2 >>
rect 2800 800 3100 810
rect 1080 780 1160 790
rect 2000 780 2080 790
rect 3820 780 3900 790
rect 4740 780 4820 790
rect 1060 700 1080 780
rect 1160 700 2000 780
rect 2080 700 2800 780
rect 3100 700 3820 780
rect 3900 700 4740 780
rect 4820 700 4840 780
rect 1080 690 1160 700
rect 2000 690 2080 700
rect 3820 690 3900 700
rect 4740 690 4820 700
rect 2800 590 3100 600
<< via2 >>
rect 2800 780 3100 800
rect 2800 700 2920 780
rect 2920 700 3000 780
rect 3000 700 3100 780
rect 2800 600 3100 700
<< metal3 >>
rect 2800 805 3100 1200
rect 2790 800 3110 805
rect 2790 600 2800 800
rect 3100 600 3110 800
rect 2790 595 3110 600
use sky130_fd_pr__nfet_01v8_lvt_J9QE6F  sky130_fd_pr__nfet_01v8_lvt_J9QE6F_1
timestamp 1672262880
transform 1 0 2726 0 1 299
box -2686 -279 2686 279
use sky130_fd_pr__nfet_01v8_lvt_M93XMJ  sky130_fd_pr__nfet_01v8_lvt_M93XMJ_0
timestamp 1672262880
transform 1 0 2726 0 1 759
box -2686 -279 2686 279
<< labels >>
flabel space 1080 -180 1180 -20 0 FreeSans 800 0 0 0 S
flabel space 1980 -160 2080 0 0 FreeSans 800 0 0 0 S
flabel space 2900 -140 3000 20 0 FreeSans 800 0 0 0 S
flabel space 3820 -140 3920 20 0 FreeSans 800 0 0 0 S
flabel space 4740 -160 4840 0 0 FreeSans 800 0 0 0 S
flabel space 1520 -180 1620 -20 0 FreeSans 800 0 0 0 D
flabel space 2440 -180 2540 -20 0 FreeSans 800 0 0 0 D
flabel space 3360 -140 3460 20 0 FreeSans 800 0 0 0 D
flabel space 4280 -120 4380 40 0 FreeSans 800 0 0 0 D
flabel space 620 -200 720 -40 0 FreeSans 800 0 0 0 D
<< end >>
