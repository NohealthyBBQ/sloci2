magic
tech sky130A
magscale 1 2
timestamp 1661879915
<< nwell >>
rect -1273 -2831 1273 2831
<< pmoslvt >>
rect -1077 1483 -977 2683
rect -919 1483 -819 2683
rect -761 1483 -661 2683
rect -603 1483 -503 2683
rect -445 1483 -345 2683
rect -287 1483 -187 2683
rect -129 1483 -29 2683
rect 29 1483 129 2683
rect 187 1483 287 2683
rect 345 1483 445 2683
rect 503 1483 603 2683
rect 661 1483 761 2683
rect 819 1483 919 2683
rect 977 1483 1077 2683
rect -1077 118 -977 1318
rect -919 118 -819 1318
rect -761 118 -661 1318
rect -603 118 -503 1318
rect -445 118 -345 1318
rect -287 118 -187 1318
rect -129 118 -29 1318
rect 29 118 129 1318
rect 187 118 287 1318
rect 345 118 445 1318
rect 503 118 603 1318
rect 661 118 761 1318
rect 819 118 919 1318
rect 977 118 1077 1318
rect -1077 -1247 -977 -47
rect -919 -1247 -819 -47
rect -761 -1247 -661 -47
rect -603 -1247 -503 -47
rect -445 -1247 -345 -47
rect -287 -1247 -187 -47
rect -129 -1247 -29 -47
rect 29 -1247 129 -47
rect 187 -1247 287 -47
rect 345 -1247 445 -47
rect 503 -1247 603 -47
rect 661 -1247 761 -47
rect 819 -1247 919 -47
rect 977 -1247 1077 -47
rect -1077 -2612 -977 -1412
rect -919 -2612 -819 -1412
rect -761 -2612 -661 -1412
rect -603 -2612 -503 -1412
rect -445 -2612 -345 -1412
rect -287 -2612 -187 -1412
rect -129 -2612 -29 -1412
rect 29 -2612 129 -1412
rect 187 -2612 287 -1412
rect 345 -2612 445 -1412
rect 503 -2612 603 -1412
rect 661 -2612 761 -1412
rect 819 -2612 919 -1412
rect 977 -2612 1077 -1412
<< pdiff >>
rect -1135 2671 -1077 2683
rect -1135 1495 -1123 2671
rect -1089 1495 -1077 2671
rect -1135 1483 -1077 1495
rect -977 2671 -919 2683
rect -977 1495 -965 2671
rect -931 1495 -919 2671
rect -977 1483 -919 1495
rect -819 2671 -761 2683
rect -819 1495 -807 2671
rect -773 1495 -761 2671
rect -819 1483 -761 1495
rect -661 2671 -603 2683
rect -661 1495 -649 2671
rect -615 1495 -603 2671
rect -661 1483 -603 1495
rect -503 2671 -445 2683
rect -503 1495 -491 2671
rect -457 1495 -445 2671
rect -503 1483 -445 1495
rect -345 2671 -287 2683
rect -345 1495 -333 2671
rect -299 1495 -287 2671
rect -345 1483 -287 1495
rect -187 2671 -129 2683
rect -187 1495 -175 2671
rect -141 1495 -129 2671
rect -187 1483 -129 1495
rect -29 2671 29 2683
rect -29 1495 -17 2671
rect 17 1495 29 2671
rect -29 1483 29 1495
rect 129 2671 187 2683
rect 129 1495 141 2671
rect 175 1495 187 2671
rect 129 1483 187 1495
rect 287 2671 345 2683
rect 287 1495 299 2671
rect 333 1495 345 2671
rect 287 1483 345 1495
rect 445 2671 503 2683
rect 445 1495 457 2671
rect 491 1495 503 2671
rect 445 1483 503 1495
rect 603 2671 661 2683
rect 603 1495 615 2671
rect 649 1495 661 2671
rect 603 1483 661 1495
rect 761 2671 819 2683
rect 761 1495 773 2671
rect 807 1495 819 2671
rect 761 1483 819 1495
rect 919 2671 977 2683
rect 919 1495 931 2671
rect 965 1495 977 2671
rect 919 1483 977 1495
rect 1077 2671 1135 2683
rect 1077 1495 1089 2671
rect 1123 1495 1135 2671
rect 1077 1483 1135 1495
rect -1135 1306 -1077 1318
rect -1135 130 -1123 1306
rect -1089 130 -1077 1306
rect -1135 118 -1077 130
rect -977 1306 -919 1318
rect -977 130 -965 1306
rect -931 130 -919 1306
rect -977 118 -919 130
rect -819 1306 -761 1318
rect -819 130 -807 1306
rect -773 130 -761 1306
rect -819 118 -761 130
rect -661 1306 -603 1318
rect -661 130 -649 1306
rect -615 130 -603 1306
rect -661 118 -603 130
rect -503 1306 -445 1318
rect -503 130 -491 1306
rect -457 130 -445 1306
rect -503 118 -445 130
rect -345 1306 -287 1318
rect -345 130 -333 1306
rect -299 130 -287 1306
rect -345 118 -287 130
rect -187 1306 -129 1318
rect -187 130 -175 1306
rect -141 130 -129 1306
rect -187 118 -129 130
rect -29 1306 29 1318
rect -29 130 -17 1306
rect 17 130 29 1306
rect -29 118 29 130
rect 129 1306 187 1318
rect 129 130 141 1306
rect 175 130 187 1306
rect 129 118 187 130
rect 287 1306 345 1318
rect 287 130 299 1306
rect 333 130 345 1306
rect 287 118 345 130
rect 445 1306 503 1318
rect 445 130 457 1306
rect 491 130 503 1306
rect 445 118 503 130
rect 603 1306 661 1318
rect 603 130 615 1306
rect 649 130 661 1306
rect 603 118 661 130
rect 761 1306 819 1318
rect 761 130 773 1306
rect 807 130 819 1306
rect 761 118 819 130
rect 919 1306 977 1318
rect 919 130 931 1306
rect 965 130 977 1306
rect 919 118 977 130
rect 1077 1306 1135 1318
rect 1077 130 1089 1306
rect 1123 130 1135 1306
rect 1077 118 1135 130
rect -1135 -59 -1077 -47
rect -1135 -1235 -1123 -59
rect -1089 -1235 -1077 -59
rect -1135 -1247 -1077 -1235
rect -977 -59 -919 -47
rect -977 -1235 -965 -59
rect -931 -1235 -919 -59
rect -977 -1247 -919 -1235
rect -819 -59 -761 -47
rect -819 -1235 -807 -59
rect -773 -1235 -761 -59
rect -819 -1247 -761 -1235
rect -661 -59 -603 -47
rect -661 -1235 -649 -59
rect -615 -1235 -603 -59
rect -661 -1247 -603 -1235
rect -503 -59 -445 -47
rect -503 -1235 -491 -59
rect -457 -1235 -445 -59
rect -503 -1247 -445 -1235
rect -345 -59 -287 -47
rect -345 -1235 -333 -59
rect -299 -1235 -287 -59
rect -345 -1247 -287 -1235
rect -187 -59 -129 -47
rect -187 -1235 -175 -59
rect -141 -1235 -129 -59
rect -187 -1247 -129 -1235
rect -29 -59 29 -47
rect -29 -1235 -17 -59
rect 17 -1235 29 -59
rect -29 -1247 29 -1235
rect 129 -59 187 -47
rect 129 -1235 141 -59
rect 175 -1235 187 -59
rect 129 -1247 187 -1235
rect 287 -59 345 -47
rect 287 -1235 299 -59
rect 333 -1235 345 -59
rect 287 -1247 345 -1235
rect 445 -59 503 -47
rect 445 -1235 457 -59
rect 491 -1235 503 -59
rect 445 -1247 503 -1235
rect 603 -59 661 -47
rect 603 -1235 615 -59
rect 649 -1235 661 -59
rect 603 -1247 661 -1235
rect 761 -59 819 -47
rect 761 -1235 773 -59
rect 807 -1235 819 -59
rect 761 -1247 819 -1235
rect 919 -59 977 -47
rect 919 -1235 931 -59
rect 965 -1235 977 -59
rect 919 -1247 977 -1235
rect 1077 -59 1135 -47
rect 1077 -1235 1089 -59
rect 1123 -1235 1135 -59
rect 1077 -1247 1135 -1235
rect -1135 -1424 -1077 -1412
rect -1135 -2600 -1123 -1424
rect -1089 -2600 -1077 -1424
rect -1135 -2612 -1077 -2600
rect -977 -1424 -919 -1412
rect -977 -2600 -965 -1424
rect -931 -2600 -919 -1424
rect -977 -2612 -919 -2600
rect -819 -1424 -761 -1412
rect -819 -2600 -807 -1424
rect -773 -2600 -761 -1424
rect -819 -2612 -761 -2600
rect -661 -1424 -603 -1412
rect -661 -2600 -649 -1424
rect -615 -2600 -603 -1424
rect -661 -2612 -603 -2600
rect -503 -1424 -445 -1412
rect -503 -2600 -491 -1424
rect -457 -2600 -445 -1424
rect -503 -2612 -445 -2600
rect -345 -1424 -287 -1412
rect -345 -2600 -333 -1424
rect -299 -2600 -287 -1424
rect -345 -2612 -287 -2600
rect -187 -1424 -129 -1412
rect -187 -2600 -175 -1424
rect -141 -2600 -129 -1424
rect -187 -2612 -129 -2600
rect -29 -1424 29 -1412
rect -29 -2600 -17 -1424
rect 17 -2600 29 -1424
rect -29 -2612 29 -2600
rect 129 -1424 187 -1412
rect 129 -2600 141 -1424
rect 175 -2600 187 -1424
rect 129 -2612 187 -2600
rect 287 -1424 345 -1412
rect 287 -2600 299 -1424
rect 333 -2600 345 -1424
rect 287 -2612 345 -2600
rect 445 -1424 503 -1412
rect 445 -2600 457 -1424
rect 491 -2600 503 -1424
rect 445 -2612 503 -2600
rect 603 -1424 661 -1412
rect 603 -2600 615 -1424
rect 649 -2600 661 -1424
rect 603 -2612 661 -2600
rect 761 -1424 819 -1412
rect 761 -2600 773 -1424
rect 807 -2600 819 -1424
rect 761 -2612 819 -2600
rect 919 -1424 977 -1412
rect 919 -2600 931 -1424
rect 965 -2600 977 -1424
rect 919 -2612 977 -2600
rect 1077 -1424 1135 -1412
rect 1077 -2600 1089 -1424
rect 1123 -2600 1135 -1424
rect 1077 -2612 1135 -2600
<< pdiffc >>
rect -1123 1495 -1089 2671
rect -965 1495 -931 2671
rect -807 1495 -773 2671
rect -649 1495 -615 2671
rect -491 1495 -457 2671
rect -333 1495 -299 2671
rect -175 1495 -141 2671
rect -17 1495 17 2671
rect 141 1495 175 2671
rect 299 1495 333 2671
rect 457 1495 491 2671
rect 615 1495 649 2671
rect 773 1495 807 2671
rect 931 1495 965 2671
rect 1089 1495 1123 2671
rect -1123 130 -1089 1306
rect -965 130 -931 1306
rect -807 130 -773 1306
rect -649 130 -615 1306
rect -491 130 -457 1306
rect -333 130 -299 1306
rect -175 130 -141 1306
rect -17 130 17 1306
rect 141 130 175 1306
rect 299 130 333 1306
rect 457 130 491 1306
rect 615 130 649 1306
rect 773 130 807 1306
rect 931 130 965 1306
rect 1089 130 1123 1306
rect -1123 -1235 -1089 -59
rect -965 -1235 -931 -59
rect -807 -1235 -773 -59
rect -649 -1235 -615 -59
rect -491 -1235 -457 -59
rect -333 -1235 -299 -59
rect -175 -1235 -141 -59
rect -17 -1235 17 -59
rect 141 -1235 175 -59
rect 299 -1235 333 -59
rect 457 -1235 491 -59
rect 615 -1235 649 -59
rect 773 -1235 807 -59
rect 931 -1235 965 -59
rect 1089 -1235 1123 -59
rect -1123 -2600 -1089 -1424
rect -965 -2600 -931 -1424
rect -807 -2600 -773 -1424
rect -649 -2600 -615 -1424
rect -491 -2600 -457 -1424
rect -333 -2600 -299 -1424
rect -175 -2600 -141 -1424
rect -17 -2600 17 -1424
rect 141 -2600 175 -1424
rect 299 -2600 333 -1424
rect 457 -2600 491 -1424
rect 615 -2600 649 -1424
rect 773 -2600 807 -1424
rect 931 -2600 965 -1424
rect 1089 -2600 1123 -1424
<< nsubdiff >>
rect -1237 2761 -1141 2795
rect 1141 2761 1237 2795
rect -1237 2699 -1203 2761
rect 1203 2699 1237 2761
rect -1237 -2761 -1203 -2699
rect 1203 -2761 1237 -2699
rect -1237 -2795 -1141 -2761
rect 1141 -2795 1237 -2761
<< nsubdiffcont >>
rect -1141 2761 1141 2795
rect -1237 -2699 -1203 2699
rect 1203 -2699 1237 2699
rect -1141 -2795 1141 -2761
<< poly >>
rect -1077 2683 -977 2709
rect -919 2683 -819 2709
rect -761 2683 -661 2709
rect -603 2683 -503 2709
rect -445 2683 -345 2709
rect -287 2683 -187 2709
rect -129 2683 -29 2709
rect 29 2683 129 2709
rect 187 2683 287 2709
rect 345 2683 445 2709
rect 503 2683 603 2709
rect 661 2683 761 2709
rect 819 2683 919 2709
rect 977 2683 1077 2709
rect -1077 1436 -977 1483
rect -1077 1402 -1061 1436
rect -993 1402 -977 1436
rect -1077 1386 -977 1402
rect -919 1436 -819 1483
rect -919 1402 -903 1436
rect -835 1402 -819 1436
rect -919 1386 -819 1402
rect -761 1436 -661 1483
rect -761 1402 -745 1436
rect -677 1402 -661 1436
rect -761 1386 -661 1402
rect -603 1436 -503 1483
rect -603 1402 -587 1436
rect -519 1402 -503 1436
rect -603 1386 -503 1402
rect -445 1436 -345 1483
rect -445 1402 -429 1436
rect -361 1402 -345 1436
rect -445 1386 -345 1402
rect -287 1436 -187 1483
rect -287 1402 -271 1436
rect -203 1402 -187 1436
rect -287 1386 -187 1402
rect -129 1436 -29 1483
rect -129 1402 -113 1436
rect -45 1402 -29 1436
rect -129 1386 -29 1402
rect 29 1436 129 1483
rect 29 1402 45 1436
rect 113 1402 129 1436
rect 29 1386 129 1402
rect 187 1436 287 1483
rect 187 1402 203 1436
rect 271 1402 287 1436
rect 187 1386 287 1402
rect 345 1436 445 1483
rect 345 1402 361 1436
rect 429 1402 445 1436
rect 345 1386 445 1402
rect 503 1436 603 1483
rect 503 1402 519 1436
rect 587 1402 603 1436
rect 503 1386 603 1402
rect 661 1436 761 1483
rect 661 1402 677 1436
rect 745 1402 761 1436
rect 661 1386 761 1402
rect 819 1436 919 1483
rect 819 1402 835 1436
rect 903 1402 919 1436
rect 819 1386 919 1402
rect 977 1436 1077 1483
rect 977 1402 993 1436
rect 1061 1402 1077 1436
rect 977 1386 1077 1402
rect -1077 1318 -977 1344
rect -919 1318 -819 1344
rect -761 1318 -661 1344
rect -603 1318 -503 1344
rect -445 1318 -345 1344
rect -287 1318 -187 1344
rect -129 1318 -29 1344
rect 29 1318 129 1344
rect 187 1318 287 1344
rect 345 1318 445 1344
rect 503 1318 603 1344
rect 661 1318 761 1344
rect 819 1318 919 1344
rect 977 1318 1077 1344
rect -1077 71 -977 118
rect -1077 37 -1061 71
rect -993 37 -977 71
rect -1077 21 -977 37
rect -919 71 -819 118
rect -919 37 -903 71
rect -835 37 -819 71
rect -919 21 -819 37
rect -761 71 -661 118
rect -761 37 -745 71
rect -677 37 -661 71
rect -761 21 -661 37
rect -603 71 -503 118
rect -603 37 -587 71
rect -519 37 -503 71
rect -603 21 -503 37
rect -445 71 -345 118
rect -445 37 -429 71
rect -361 37 -345 71
rect -445 21 -345 37
rect -287 71 -187 118
rect -287 37 -271 71
rect -203 37 -187 71
rect -287 21 -187 37
rect -129 71 -29 118
rect -129 37 -113 71
rect -45 37 -29 71
rect -129 21 -29 37
rect 29 71 129 118
rect 29 37 45 71
rect 113 37 129 71
rect 29 21 129 37
rect 187 71 287 118
rect 187 37 203 71
rect 271 37 287 71
rect 187 21 287 37
rect 345 71 445 118
rect 345 37 361 71
rect 429 37 445 71
rect 345 21 445 37
rect 503 71 603 118
rect 503 37 519 71
rect 587 37 603 71
rect 503 21 603 37
rect 661 71 761 118
rect 661 37 677 71
rect 745 37 761 71
rect 661 21 761 37
rect 819 71 919 118
rect 819 37 835 71
rect 903 37 919 71
rect 819 21 919 37
rect 977 71 1077 118
rect 977 37 993 71
rect 1061 37 1077 71
rect 977 21 1077 37
rect -1077 -47 -977 -21
rect -919 -47 -819 -21
rect -761 -47 -661 -21
rect -603 -47 -503 -21
rect -445 -47 -345 -21
rect -287 -47 -187 -21
rect -129 -47 -29 -21
rect 29 -47 129 -21
rect 187 -47 287 -21
rect 345 -47 445 -21
rect 503 -47 603 -21
rect 661 -47 761 -21
rect 819 -47 919 -21
rect 977 -47 1077 -21
rect -1077 -1294 -977 -1247
rect -1077 -1328 -1061 -1294
rect -993 -1328 -977 -1294
rect -1077 -1344 -977 -1328
rect -919 -1294 -819 -1247
rect -919 -1328 -903 -1294
rect -835 -1328 -819 -1294
rect -919 -1344 -819 -1328
rect -761 -1294 -661 -1247
rect -761 -1328 -745 -1294
rect -677 -1328 -661 -1294
rect -761 -1344 -661 -1328
rect -603 -1294 -503 -1247
rect -603 -1328 -587 -1294
rect -519 -1328 -503 -1294
rect -603 -1344 -503 -1328
rect -445 -1294 -345 -1247
rect -445 -1328 -429 -1294
rect -361 -1328 -345 -1294
rect -445 -1344 -345 -1328
rect -287 -1294 -187 -1247
rect -287 -1328 -271 -1294
rect -203 -1328 -187 -1294
rect -287 -1344 -187 -1328
rect -129 -1294 -29 -1247
rect -129 -1328 -113 -1294
rect -45 -1328 -29 -1294
rect -129 -1344 -29 -1328
rect 29 -1294 129 -1247
rect 29 -1328 45 -1294
rect 113 -1328 129 -1294
rect 29 -1344 129 -1328
rect 187 -1294 287 -1247
rect 187 -1328 203 -1294
rect 271 -1328 287 -1294
rect 187 -1344 287 -1328
rect 345 -1294 445 -1247
rect 345 -1328 361 -1294
rect 429 -1328 445 -1294
rect 345 -1344 445 -1328
rect 503 -1294 603 -1247
rect 503 -1328 519 -1294
rect 587 -1328 603 -1294
rect 503 -1344 603 -1328
rect 661 -1294 761 -1247
rect 661 -1328 677 -1294
rect 745 -1328 761 -1294
rect 661 -1344 761 -1328
rect 819 -1294 919 -1247
rect 819 -1328 835 -1294
rect 903 -1328 919 -1294
rect 819 -1344 919 -1328
rect 977 -1294 1077 -1247
rect 977 -1328 993 -1294
rect 1061 -1328 1077 -1294
rect 977 -1344 1077 -1328
rect -1077 -1412 -977 -1386
rect -919 -1412 -819 -1386
rect -761 -1412 -661 -1386
rect -603 -1412 -503 -1386
rect -445 -1412 -345 -1386
rect -287 -1412 -187 -1386
rect -129 -1412 -29 -1386
rect 29 -1412 129 -1386
rect 187 -1412 287 -1386
rect 345 -1412 445 -1386
rect 503 -1412 603 -1386
rect 661 -1412 761 -1386
rect 819 -1412 919 -1386
rect 977 -1412 1077 -1386
rect -1077 -2659 -977 -2612
rect -1077 -2693 -1061 -2659
rect -993 -2693 -977 -2659
rect -1077 -2709 -977 -2693
rect -919 -2659 -819 -2612
rect -919 -2693 -903 -2659
rect -835 -2693 -819 -2659
rect -919 -2709 -819 -2693
rect -761 -2659 -661 -2612
rect -761 -2693 -745 -2659
rect -677 -2693 -661 -2659
rect -761 -2709 -661 -2693
rect -603 -2659 -503 -2612
rect -603 -2693 -587 -2659
rect -519 -2693 -503 -2659
rect -603 -2709 -503 -2693
rect -445 -2659 -345 -2612
rect -445 -2693 -429 -2659
rect -361 -2693 -345 -2659
rect -445 -2709 -345 -2693
rect -287 -2659 -187 -2612
rect -287 -2693 -271 -2659
rect -203 -2693 -187 -2659
rect -287 -2709 -187 -2693
rect -129 -2659 -29 -2612
rect -129 -2693 -113 -2659
rect -45 -2693 -29 -2659
rect -129 -2709 -29 -2693
rect 29 -2659 129 -2612
rect 29 -2693 45 -2659
rect 113 -2693 129 -2659
rect 29 -2709 129 -2693
rect 187 -2659 287 -2612
rect 187 -2693 203 -2659
rect 271 -2693 287 -2659
rect 187 -2709 287 -2693
rect 345 -2659 445 -2612
rect 345 -2693 361 -2659
rect 429 -2693 445 -2659
rect 345 -2709 445 -2693
rect 503 -2659 603 -2612
rect 503 -2693 519 -2659
rect 587 -2693 603 -2659
rect 503 -2709 603 -2693
rect 661 -2659 761 -2612
rect 661 -2693 677 -2659
rect 745 -2693 761 -2659
rect 661 -2709 761 -2693
rect 819 -2659 919 -2612
rect 819 -2693 835 -2659
rect 903 -2693 919 -2659
rect 819 -2709 919 -2693
rect 977 -2659 1077 -2612
rect 977 -2693 993 -2659
rect 1061 -2693 1077 -2659
rect 977 -2709 1077 -2693
<< polycont >>
rect -1061 1402 -993 1436
rect -903 1402 -835 1436
rect -745 1402 -677 1436
rect -587 1402 -519 1436
rect -429 1402 -361 1436
rect -271 1402 -203 1436
rect -113 1402 -45 1436
rect 45 1402 113 1436
rect 203 1402 271 1436
rect 361 1402 429 1436
rect 519 1402 587 1436
rect 677 1402 745 1436
rect 835 1402 903 1436
rect 993 1402 1061 1436
rect -1061 37 -993 71
rect -903 37 -835 71
rect -745 37 -677 71
rect -587 37 -519 71
rect -429 37 -361 71
rect -271 37 -203 71
rect -113 37 -45 71
rect 45 37 113 71
rect 203 37 271 71
rect 361 37 429 71
rect 519 37 587 71
rect 677 37 745 71
rect 835 37 903 71
rect 993 37 1061 71
rect -1061 -1328 -993 -1294
rect -903 -1328 -835 -1294
rect -745 -1328 -677 -1294
rect -587 -1328 -519 -1294
rect -429 -1328 -361 -1294
rect -271 -1328 -203 -1294
rect -113 -1328 -45 -1294
rect 45 -1328 113 -1294
rect 203 -1328 271 -1294
rect 361 -1328 429 -1294
rect 519 -1328 587 -1294
rect 677 -1328 745 -1294
rect 835 -1328 903 -1294
rect 993 -1328 1061 -1294
rect -1061 -2693 -993 -2659
rect -903 -2693 -835 -2659
rect -745 -2693 -677 -2659
rect -587 -2693 -519 -2659
rect -429 -2693 -361 -2659
rect -271 -2693 -203 -2659
rect -113 -2693 -45 -2659
rect 45 -2693 113 -2659
rect 203 -2693 271 -2659
rect 361 -2693 429 -2659
rect 519 -2693 587 -2659
rect 677 -2693 745 -2659
rect 835 -2693 903 -2659
rect 993 -2693 1061 -2659
<< locali >>
rect -1237 2761 -1141 2795
rect 1141 2761 1237 2795
rect -1237 2699 -1203 2761
rect 1203 2699 1237 2761
rect -1123 2671 -1089 2687
rect -1123 1479 -1089 1495
rect -965 2671 -931 2687
rect -965 1479 -931 1495
rect -807 2671 -773 2687
rect -807 1479 -773 1495
rect -649 2671 -615 2687
rect -649 1479 -615 1495
rect -491 2671 -457 2687
rect -491 1479 -457 1495
rect -333 2671 -299 2687
rect -333 1479 -299 1495
rect -175 2671 -141 2687
rect -175 1479 -141 1495
rect -17 2671 17 2687
rect -17 1479 17 1495
rect 141 2671 175 2687
rect 141 1479 175 1495
rect 299 2671 333 2687
rect 299 1479 333 1495
rect 457 2671 491 2687
rect 457 1479 491 1495
rect 615 2671 649 2687
rect 615 1479 649 1495
rect 773 2671 807 2687
rect 773 1479 807 1495
rect 931 2671 965 2687
rect 931 1479 965 1495
rect 1089 2671 1123 2687
rect 1089 1479 1123 1495
rect -1077 1402 -1061 1436
rect -993 1402 -977 1436
rect -919 1402 -903 1436
rect -835 1402 -819 1436
rect -761 1402 -745 1436
rect -677 1402 -661 1436
rect -603 1402 -587 1436
rect -519 1402 -503 1436
rect -445 1402 -429 1436
rect -361 1402 -345 1436
rect -287 1402 -271 1436
rect -203 1402 -187 1436
rect -129 1402 -113 1436
rect -45 1402 -29 1436
rect 29 1402 45 1436
rect 113 1402 129 1436
rect 187 1402 203 1436
rect 271 1402 287 1436
rect 345 1402 361 1436
rect 429 1402 445 1436
rect 503 1402 519 1436
rect 587 1402 603 1436
rect 661 1402 677 1436
rect 745 1402 761 1436
rect 819 1402 835 1436
rect 903 1402 919 1436
rect 977 1402 993 1436
rect 1061 1402 1077 1436
rect -1123 1306 -1089 1322
rect -1123 114 -1089 130
rect -965 1306 -931 1322
rect -965 114 -931 130
rect -807 1306 -773 1322
rect -807 114 -773 130
rect -649 1306 -615 1322
rect -649 114 -615 130
rect -491 1306 -457 1322
rect -491 114 -457 130
rect -333 1306 -299 1322
rect -333 114 -299 130
rect -175 1306 -141 1322
rect -175 114 -141 130
rect -17 1306 17 1322
rect -17 114 17 130
rect 141 1306 175 1322
rect 141 114 175 130
rect 299 1306 333 1322
rect 299 114 333 130
rect 457 1306 491 1322
rect 457 114 491 130
rect 615 1306 649 1322
rect 615 114 649 130
rect 773 1306 807 1322
rect 773 114 807 130
rect 931 1306 965 1322
rect 931 114 965 130
rect 1089 1306 1123 1322
rect 1089 114 1123 130
rect -1077 37 -1061 71
rect -993 37 -977 71
rect -919 37 -903 71
rect -835 37 -819 71
rect -761 37 -745 71
rect -677 37 -661 71
rect -603 37 -587 71
rect -519 37 -503 71
rect -445 37 -429 71
rect -361 37 -345 71
rect -287 37 -271 71
rect -203 37 -187 71
rect -129 37 -113 71
rect -45 37 -29 71
rect 29 37 45 71
rect 113 37 129 71
rect 187 37 203 71
rect 271 37 287 71
rect 345 37 361 71
rect 429 37 445 71
rect 503 37 519 71
rect 587 37 603 71
rect 661 37 677 71
rect 745 37 761 71
rect 819 37 835 71
rect 903 37 919 71
rect 977 37 993 71
rect 1061 37 1077 71
rect -1123 -59 -1089 -43
rect -1123 -1251 -1089 -1235
rect -965 -59 -931 -43
rect -965 -1251 -931 -1235
rect -807 -59 -773 -43
rect -807 -1251 -773 -1235
rect -649 -59 -615 -43
rect -649 -1251 -615 -1235
rect -491 -59 -457 -43
rect -491 -1251 -457 -1235
rect -333 -59 -299 -43
rect -333 -1251 -299 -1235
rect -175 -59 -141 -43
rect -175 -1251 -141 -1235
rect -17 -59 17 -43
rect -17 -1251 17 -1235
rect 141 -59 175 -43
rect 141 -1251 175 -1235
rect 299 -59 333 -43
rect 299 -1251 333 -1235
rect 457 -59 491 -43
rect 457 -1251 491 -1235
rect 615 -59 649 -43
rect 615 -1251 649 -1235
rect 773 -59 807 -43
rect 773 -1251 807 -1235
rect 931 -59 965 -43
rect 931 -1251 965 -1235
rect 1089 -59 1123 -43
rect 1089 -1251 1123 -1235
rect -1077 -1328 -1061 -1294
rect -993 -1328 -977 -1294
rect -919 -1328 -903 -1294
rect -835 -1328 -819 -1294
rect -761 -1328 -745 -1294
rect -677 -1328 -661 -1294
rect -603 -1328 -587 -1294
rect -519 -1328 -503 -1294
rect -445 -1328 -429 -1294
rect -361 -1328 -345 -1294
rect -287 -1328 -271 -1294
rect -203 -1328 -187 -1294
rect -129 -1328 -113 -1294
rect -45 -1328 -29 -1294
rect 29 -1328 45 -1294
rect 113 -1328 129 -1294
rect 187 -1328 203 -1294
rect 271 -1328 287 -1294
rect 345 -1328 361 -1294
rect 429 -1328 445 -1294
rect 503 -1328 519 -1294
rect 587 -1328 603 -1294
rect 661 -1328 677 -1294
rect 745 -1328 761 -1294
rect 819 -1328 835 -1294
rect 903 -1328 919 -1294
rect 977 -1328 993 -1294
rect 1061 -1328 1077 -1294
rect -1123 -1424 -1089 -1408
rect -1123 -2616 -1089 -2600
rect -965 -1424 -931 -1408
rect -965 -2616 -931 -2600
rect -807 -1424 -773 -1408
rect -807 -2616 -773 -2600
rect -649 -1424 -615 -1408
rect -649 -2616 -615 -2600
rect -491 -1424 -457 -1408
rect -491 -2616 -457 -2600
rect -333 -1424 -299 -1408
rect -333 -2616 -299 -2600
rect -175 -1424 -141 -1408
rect -175 -2616 -141 -2600
rect -17 -1424 17 -1408
rect -17 -2616 17 -2600
rect 141 -1424 175 -1408
rect 141 -2616 175 -2600
rect 299 -1424 333 -1408
rect 299 -2616 333 -2600
rect 457 -1424 491 -1408
rect 457 -2616 491 -2600
rect 615 -1424 649 -1408
rect 615 -2616 649 -2600
rect 773 -1424 807 -1408
rect 773 -2616 807 -2600
rect 931 -1424 965 -1408
rect 931 -2616 965 -2600
rect 1089 -1424 1123 -1408
rect 1089 -2616 1123 -2600
rect -1077 -2693 -1061 -2659
rect -993 -2693 -977 -2659
rect -919 -2693 -903 -2659
rect -835 -2693 -819 -2659
rect -761 -2693 -745 -2659
rect -677 -2693 -661 -2659
rect -603 -2693 -587 -2659
rect -519 -2693 -503 -2659
rect -445 -2693 -429 -2659
rect -361 -2693 -345 -2659
rect -287 -2693 -271 -2659
rect -203 -2693 -187 -2659
rect -129 -2693 -113 -2659
rect -45 -2693 -29 -2659
rect 29 -2693 45 -2659
rect 113 -2693 129 -2659
rect 187 -2693 203 -2659
rect 271 -2693 287 -2659
rect 345 -2693 361 -2659
rect 429 -2693 445 -2659
rect 503 -2693 519 -2659
rect 587 -2693 603 -2659
rect 661 -2693 677 -2659
rect 745 -2693 761 -2659
rect 819 -2693 835 -2659
rect 903 -2693 919 -2659
rect 977 -2693 993 -2659
rect 1061 -2693 1077 -2659
rect -1237 -2761 -1203 -2699
rect 1203 -2761 1237 -2699
rect -1237 -2795 -1141 -2761
rect 1141 -2795 1237 -2761
<< viali >>
rect -1123 1495 -1089 2671
rect -965 1495 -931 2671
rect -807 1495 -773 2671
rect -649 1495 -615 2671
rect -491 1495 -457 2671
rect -333 1495 -299 2671
rect -175 1495 -141 2671
rect -17 1495 17 2671
rect 141 1495 175 2671
rect 299 1495 333 2671
rect 457 1495 491 2671
rect 615 1495 649 2671
rect 773 1495 807 2671
rect 931 1495 965 2671
rect 1089 1495 1123 2671
rect -1061 1402 -993 1436
rect -903 1402 -835 1436
rect -745 1402 -677 1436
rect -587 1402 -519 1436
rect -429 1402 -361 1436
rect -271 1402 -203 1436
rect -113 1402 -45 1436
rect 45 1402 113 1436
rect 203 1402 271 1436
rect 361 1402 429 1436
rect 519 1402 587 1436
rect 677 1402 745 1436
rect 835 1402 903 1436
rect 993 1402 1061 1436
rect -1123 130 -1089 1306
rect -965 130 -931 1306
rect -807 130 -773 1306
rect -649 130 -615 1306
rect -491 130 -457 1306
rect -333 130 -299 1306
rect -175 130 -141 1306
rect -17 130 17 1306
rect 141 130 175 1306
rect 299 130 333 1306
rect 457 130 491 1306
rect 615 130 649 1306
rect 773 130 807 1306
rect 931 130 965 1306
rect 1089 130 1123 1306
rect -1061 37 -993 71
rect -903 37 -835 71
rect -745 37 -677 71
rect -587 37 -519 71
rect -429 37 -361 71
rect -271 37 -203 71
rect -113 37 -45 71
rect 45 37 113 71
rect 203 37 271 71
rect 361 37 429 71
rect 519 37 587 71
rect 677 37 745 71
rect 835 37 903 71
rect 993 37 1061 71
rect -1123 -1235 -1089 -59
rect -965 -1235 -931 -59
rect -807 -1235 -773 -59
rect -649 -1235 -615 -59
rect -491 -1235 -457 -59
rect -333 -1235 -299 -59
rect -175 -1235 -141 -59
rect -17 -1235 17 -59
rect 141 -1235 175 -59
rect 299 -1235 333 -59
rect 457 -1235 491 -59
rect 615 -1235 649 -59
rect 773 -1235 807 -59
rect 931 -1235 965 -59
rect 1089 -1235 1123 -59
rect -1061 -1328 -993 -1294
rect -903 -1328 -835 -1294
rect -745 -1328 -677 -1294
rect -587 -1328 -519 -1294
rect -429 -1328 -361 -1294
rect -271 -1328 -203 -1294
rect -113 -1328 -45 -1294
rect 45 -1328 113 -1294
rect 203 -1328 271 -1294
rect 361 -1328 429 -1294
rect 519 -1328 587 -1294
rect 677 -1328 745 -1294
rect 835 -1328 903 -1294
rect 993 -1328 1061 -1294
rect -1123 -2600 -1089 -1424
rect -965 -2600 -931 -1424
rect -807 -2600 -773 -1424
rect -649 -2600 -615 -1424
rect -491 -2600 -457 -1424
rect -333 -2600 -299 -1424
rect -175 -2600 -141 -1424
rect -17 -2600 17 -1424
rect 141 -2600 175 -1424
rect 299 -2600 333 -1424
rect 457 -2600 491 -1424
rect 615 -2600 649 -1424
rect 773 -2600 807 -1424
rect 931 -2600 965 -1424
rect 1089 -2600 1123 -1424
rect -1061 -2693 -993 -2659
rect -903 -2693 -835 -2659
rect -745 -2693 -677 -2659
rect -587 -2693 -519 -2659
rect -429 -2693 -361 -2659
rect -271 -2693 -203 -2659
rect -113 -2693 -45 -2659
rect 45 -2693 113 -2659
rect 203 -2693 271 -2659
rect 361 -2693 429 -2659
rect 519 -2693 587 -2659
rect 677 -2693 745 -2659
rect 835 -2693 903 -2659
rect 993 -2693 1061 -2659
<< metal1 >>
rect -1129 2671 -1083 2683
rect -1129 1495 -1123 2671
rect -1089 1495 -1083 2671
rect -1129 1483 -1083 1495
rect -971 2671 -925 2683
rect -971 1495 -965 2671
rect -931 1495 -925 2671
rect -971 1483 -925 1495
rect -813 2671 -767 2683
rect -813 1495 -807 2671
rect -773 1495 -767 2671
rect -813 1483 -767 1495
rect -655 2671 -609 2683
rect -655 1495 -649 2671
rect -615 1495 -609 2671
rect -655 1483 -609 1495
rect -497 2671 -451 2683
rect -497 1495 -491 2671
rect -457 1495 -451 2671
rect -497 1483 -451 1495
rect -339 2671 -293 2683
rect -339 1495 -333 2671
rect -299 1495 -293 2671
rect -339 1483 -293 1495
rect -181 2671 -135 2683
rect -181 1495 -175 2671
rect -141 1495 -135 2671
rect -181 1483 -135 1495
rect -23 2671 23 2683
rect -23 1495 -17 2671
rect 17 1495 23 2671
rect -23 1483 23 1495
rect 135 2671 181 2683
rect 135 1495 141 2671
rect 175 1495 181 2671
rect 135 1483 181 1495
rect 293 2671 339 2683
rect 293 1495 299 2671
rect 333 1495 339 2671
rect 293 1483 339 1495
rect 451 2671 497 2683
rect 451 1495 457 2671
rect 491 1495 497 2671
rect 451 1483 497 1495
rect 609 2671 655 2683
rect 609 1495 615 2671
rect 649 1495 655 2671
rect 609 1483 655 1495
rect 767 2671 813 2683
rect 767 1495 773 2671
rect 807 1495 813 2671
rect 767 1483 813 1495
rect 925 2671 971 2683
rect 925 1495 931 2671
rect 965 1495 971 2671
rect 925 1483 971 1495
rect 1083 2671 1129 2683
rect 1083 1495 1089 2671
rect 1123 1495 1129 2671
rect 1083 1483 1129 1495
rect -1073 1436 -981 1442
rect -1073 1402 -1061 1436
rect -993 1402 -981 1436
rect -1073 1396 -981 1402
rect -915 1436 -823 1442
rect -915 1402 -903 1436
rect -835 1402 -823 1436
rect -915 1396 -823 1402
rect -757 1436 -665 1442
rect -757 1402 -745 1436
rect -677 1402 -665 1436
rect -757 1396 -665 1402
rect -599 1436 -507 1442
rect -599 1402 -587 1436
rect -519 1402 -507 1436
rect -599 1396 -507 1402
rect -441 1436 -349 1442
rect -441 1402 -429 1436
rect -361 1402 -349 1436
rect -441 1396 -349 1402
rect -283 1436 -191 1442
rect -283 1402 -271 1436
rect -203 1402 -191 1436
rect -283 1396 -191 1402
rect -125 1436 -33 1442
rect -125 1402 -113 1436
rect -45 1402 -33 1436
rect -125 1396 -33 1402
rect 33 1436 125 1442
rect 33 1402 45 1436
rect 113 1402 125 1436
rect 33 1396 125 1402
rect 191 1436 283 1442
rect 191 1402 203 1436
rect 271 1402 283 1436
rect 191 1396 283 1402
rect 349 1436 441 1442
rect 349 1402 361 1436
rect 429 1402 441 1436
rect 349 1396 441 1402
rect 507 1436 599 1442
rect 507 1402 519 1436
rect 587 1402 599 1436
rect 507 1396 599 1402
rect 665 1436 757 1442
rect 665 1402 677 1436
rect 745 1402 757 1436
rect 665 1396 757 1402
rect 823 1436 915 1442
rect 823 1402 835 1436
rect 903 1402 915 1436
rect 823 1396 915 1402
rect 981 1436 1073 1442
rect 981 1402 993 1436
rect 1061 1402 1073 1436
rect 981 1396 1073 1402
rect -1129 1306 -1083 1318
rect -1129 130 -1123 1306
rect -1089 130 -1083 1306
rect -1129 118 -1083 130
rect -971 1306 -925 1318
rect -971 130 -965 1306
rect -931 130 -925 1306
rect -971 118 -925 130
rect -813 1306 -767 1318
rect -813 130 -807 1306
rect -773 130 -767 1306
rect -813 118 -767 130
rect -655 1306 -609 1318
rect -655 130 -649 1306
rect -615 130 -609 1306
rect -655 118 -609 130
rect -497 1306 -451 1318
rect -497 130 -491 1306
rect -457 130 -451 1306
rect -497 118 -451 130
rect -339 1306 -293 1318
rect -339 130 -333 1306
rect -299 130 -293 1306
rect -339 118 -293 130
rect -181 1306 -135 1318
rect -181 130 -175 1306
rect -141 130 -135 1306
rect -181 118 -135 130
rect -23 1306 23 1318
rect -23 130 -17 1306
rect 17 130 23 1306
rect -23 118 23 130
rect 135 1306 181 1318
rect 135 130 141 1306
rect 175 130 181 1306
rect 135 118 181 130
rect 293 1306 339 1318
rect 293 130 299 1306
rect 333 130 339 1306
rect 293 118 339 130
rect 451 1306 497 1318
rect 451 130 457 1306
rect 491 130 497 1306
rect 451 118 497 130
rect 609 1306 655 1318
rect 609 130 615 1306
rect 649 130 655 1306
rect 609 118 655 130
rect 767 1306 813 1318
rect 767 130 773 1306
rect 807 130 813 1306
rect 767 118 813 130
rect 925 1306 971 1318
rect 925 130 931 1306
rect 965 130 971 1306
rect 925 118 971 130
rect 1083 1306 1129 1318
rect 1083 130 1089 1306
rect 1123 130 1129 1306
rect 1083 118 1129 130
rect -1073 71 -981 77
rect -1073 37 -1061 71
rect -993 37 -981 71
rect -1073 31 -981 37
rect -915 71 -823 77
rect -915 37 -903 71
rect -835 37 -823 71
rect -915 31 -823 37
rect -757 71 -665 77
rect -757 37 -745 71
rect -677 37 -665 71
rect -757 31 -665 37
rect -599 71 -507 77
rect -599 37 -587 71
rect -519 37 -507 71
rect -599 31 -507 37
rect -441 71 -349 77
rect -441 37 -429 71
rect -361 37 -349 71
rect -441 31 -349 37
rect -283 71 -191 77
rect -283 37 -271 71
rect -203 37 -191 71
rect -283 31 -191 37
rect -125 71 -33 77
rect -125 37 -113 71
rect -45 37 -33 71
rect -125 31 -33 37
rect 33 71 125 77
rect 33 37 45 71
rect 113 37 125 71
rect 33 31 125 37
rect 191 71 283 77
rect 191 37 203 71
rect 271 37 283 71
rect 191 31 283 37
rect 349 71 441 77
rect 349 37 361 71
rect 429 37 441 71
rect 349 31 441 37
rect 507 71 599 77
rect 507 37 519 71
rect 587 37 599 71
rect 507 31 599 37
rect 665 71 757 77
rect 665 37 677 71
rect 745 37 757 71
rect 665 31 757 37
rect 823 71 915 77
rect 823 37 835 71
rect 903 37 915 71
rect 823 31 915 37
rect 981 71 1073 77
rect 981 37 993 71
rect 1061 37 1073 71
rect 981 31 1073 37
rect -1129 -59 -1083 -47
rect -1129 -1235 -1123 -59
rect -1089 -1235 -1083 -59
rect -1129 -1247 -1083 -1235
rect -971 -59 -925 -47
rect -971 -1235 -965 -59
rect -931 -1235 -925 -59
rect -971 -1247 -925 -1235
rect -813 -59 -767 -47
rect -813 -1235 -807 -59
rect -773 -1235 -767 -59
rect -813 -1247 -767 -1235
rect -655 -59 -609 -47
rect -655 -1235 -649 -59
rect -615 -1235 -609 -59
rect -655 -1247 -609 -1235
rect -497 -59 -451 -47
rect -497 -1235 -491 -59
rect -457 -1235 -451 -59
rect -497 -1247 -451 -1235
rect -339 -59 -293 -47
rect -339 -1235 -333 -59
rect -299 -1235 -293 -59
rect -339 -1247 -293 -1235
rect -181 -59 -135 -47
rect -181 -1235 -175 -59
rect -141 -1235 -135 -59
rect -181 -1247 -135 -1235
rect -23 -59 23 -47
rect -23 -1235 -17 -59
rect 17 -1235 23 -59
rect -23 -1247 23 -1235
rect 135 -59 181 -47
rect 135 -1235 141 -59
rect 175 -1235 181 -59
rect 135 -1247 181 -1235
rect 293 -59 339 -47
rect 293 -1235 299 -59
rect 333 -1235 339 -59
rect 293 -1247 339 -1235
rect 451 -59 497 -47
rect 451 -1235 457 -59
rect 491 -1235 497 -59
rect 451 -1247 497 -1235
rect 609 -59 655 -47
rect 609 -1235 615 -59
rect 649 -1235 655 -59
rect 609 -1247 655 -1235
rect 767 -59 813 -47
rect 767 -1235 773 -59
rect 807 -1235 813 -59
rect 767 -1247 813 -1235
rect 925 -59 971 -47
rect 925 -1235 931 -59
rect 965 -1235 971 -59
rect 925 -1247 971 -1235
rect 1083 -59 1129 -47
rect 1083 -1235 1089 -59
rect 1123 -1235 1129 -59
rect 1083 -1247 1129 -1235
rect -1073 -1294 -981 -1288
rect -1073 -1328 -1061 -1294
rect -993 -1328 -981 -1294
rect -1073 -1334 -981 -1328
rect -915 -1294 -823 -1288
rect -915 -1328 -903 -1294
rect -835 -1328 -823 -1294
rect -915 -1334 -823 -1328
rect -757 -1294 -665 -1288
rect -757 -1328 -745 -1294
rect -677 -1328 -665 -1294
rect -757 -1334 -665 -1328
rect -599 -1294 -507 -1288
rect -599 -1328 -587 -1294
rect -519 -1328 -507 -1294
rect -599 -1334 -507 -1328
rect -441 -1294 -349 -1288
rect -441 -1328 -429 -1294
rect -361 -1328 -349 -1294
rect -441 -1334 -349 -1328
rect -283 -1294 -191 -1288
rect -283 -1328 -271 -1294
rect -203 -1328 -191 -1294
rect -283 -1334 -191 -1328
rect -125 -1294 -33 -1288
rect -125 -1328 -113 -1294
rect -45 -1328 -33 -1294
rect -125 -1334 -33 -1328
rect 33 -1294 125 -1288
rect 33 -1328 45 -1294
rect 113 -1328 125 -1294
rect 33 -1334 125 -1328
rect 191 -1294 283 -1288
rect 191 -1328 203 -1294
rect 271 -1328 283 -1294
rect 191 -1334 283 -1328
rect 349 -1294 441 -1288
rect 349 -1328 361 -1294
rect 429 -1328 441 -1294
rect 349 -1334 441 -1328
rect 507 -1294 599 -1288
rect 507 -1328 519 -1294
rect 587 -1328 599 -1294
rect 507 -1334 599 -1328
rect 665 -1294 757 -1288
rect 665 -1328 677 -1294
rect 745 -1328 757 -1294
rect 665 -1334 757 -1328
rect 823 -1294 915 -1288
rect 823 -1328 835 -1294
rect 903 -1328 915 -1294
rect 823 -1334 915 -1328
rect 981 -1294 1073 -1288
rect 981 -1328 993 -1294
rect 1061 -1328 1073 -1294
rect 981 -1334 1073 -1328
rect -1129 -1424 -1083 -1412
rect -1129 -2600 -1123 -1424
rect -1089 -2600 -1083 -1424
rect -1129 -2612 -1083 -2600
rect -971 -1424 -925 -1412
rect -971 -2600 -965 -1424
rect -931 -2600 -925 -1424
rect -971 -2612 -925 -2600
rect -813 -1424 -767 -1412
rect -813 -2600 -807 -1424
rect -773 -2600 -767 -1424
rect -813 -2612 -767 -2600
rect -655 -1424 -609 -1412
rect -655 -2600 -649 -1424
rect -615 -2600 -609 -1424
rect -655 -2612 -609 -2600
rect -497 -1424 -451 -1412
rect -497 -2600 -491 -1424
rect -457 -2600 -451 -1424
rect -497 -2612 -451 -2600
rect -339 -1424 -293 -1412
rect -339 -2600 -333 -1424
rect -299 -2600 -293 -1424
rect -339 -2612 -293 -2600
rect -181 -1424 -135 -1412
rect -181 -2600 -175 -1424
rect -141 -2600 -135 -1424
rect -181 -2612 -135 -2600
rect -23 -1424 23 -1412
rect -23 -2600 -17 -1424
rect 17 -2600 23 -1424
rect -23 -2612 23 -2600
rect 135 -1424 181 -1412
rect 135 -2600 141 -1424
rect 175 -2600 181 -1424
rect 135 -2612 181 -2600
rect 293 -1424 339 -1412
rect 293 -2600 299 -1424
rect 333 -2600 339 -1424
rect 293 -2612 339 -2600
rect 451 -1424 497 -1412
rect 451 -2600 457 -1424
rect 491 -2600 497 -1424
rect 451 -2612 497 -2600
rect 609 -1424 655 -1412
rect 609 -2600 615 -1424
rect 649 -2600 655 -1424
rect 609 -2612 655 -2600
rect 767 -1424 813 -1412
rect 767 -2600 773 -1424
rect 807 -2600 813 -1424
rect 767 -2612 813 -2600
rect 925 -1424 971 -1412
rect 925 -2600 931 -1424
rect 965 -2600 971 -1424
rect 925 -2612 971 -2600
rect 1083 -1424 1129 -1412
rect 1083 -2600 1089 -1424
rect 1123 -2600 1129 -1424
rect 1083 -2612 1129 -2600
rect -1073 -2659 -981 -2653
rect -1073 -2693 -1061 -2659
rect -993 -2693 -981 -2659
rect -1073 -2699 -981 -2693
rect -915 -2659 -823 -2653
rect -915 -2693 -903 -2659
rect -835 -2693 -823 -2659
rect -915 -2699 -823 -2693
rect -757 -2659 -665 -2653
rect -757 -2693 -745 -2659
rect -677 -2693 -665 -2659
rect -757 -2699 -665 -2693
rect -599 -2659 -507 -2653
rect -599 -2693 -587 -2659
rect -519 -2693 -507 -2659
rect -599 -2699 -507 -2693
rect -441 -2659 -349 -2653
rect -441 -2693 -429 -2659
rect -361 -2693 -349 -2659
rect -441 -2699 -349 -2693
rect -283 -2659 -191 -2653
rect -283 -2693 -271 -2659
rect -203 -2693 -191 -2659
rect -283 -2699 -191 -2693
rect -125 -2659 -33 -2653
rect -125 -2693 -113 -2659
rect -45 -2693 -33 -2659
rect -125 -2699 -33 -2693
rect 33 -2659 125 -2653
rect 33 -2693 45 -2659
rect 113 -2693 125 -2659
rect 33 -2699 125 -2693
rect 191 -2659 283 -2653
rect 191 -2693 203 -2659
rect 271 -2693 283 -2659
rect 191 -2699 283 -2693
rect 349 -2659 441 -2653
rect 349 -2693 361 -2659
rect 429 -2693 441 -2659
rect 349 -2699 441 -2693
rect 507 -2659 599 -2653
rect 507 -2693 519 -2659
rect 587 -2693 599 -2659
rect 507 -2699 599 -2693
rect 665 -2659 757 -2653
rect 665 -2693 677 -2659
rect 745 -2693 757 -2659
rect 665 -2699 757 -2693
rect 823 -2659 915 -2653
rect 823 -2693 835 -2659
rect 903 -2693 915 -2659
rect 823 -2699 915 -2693
rect 981 -2659 1073 -2653
rect 981 -2693 993 -2659
rect 1061 -2693 1073 -2659
rect 981 -2699 1073 -2693
<< properties >>
string FIXED_BBOX -1220 -2778 1220 2778
string gencell sky130_fd_pr__pfet_01v8_lvt
string library sky130
string parameters w 6 l 0.5 m 4 nf 14 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 0 botc 1 poverlap 0 doverlap 1 lmin 0.35 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
