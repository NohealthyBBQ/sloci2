magic
tech sky130A
magscale 1 2
timestamp 1662690363
<< error_p >>
rect -159 372 -97 378
rect -31 372 31 378
rect 97 372 159 378
rect -159 338 -147 372
rect -31 338 -19 372
rect 97 338 109 372
rect -159 332 -97 338
rect -31 332 31 338
rect 97 332 159 338
rect -159 -338 -97 -332
rect -31 -338 31 -332
rect 97 -338 159 -332
rect -159 -372 -147 -338
rect -31 -372 -19 -338
rect 97 -372 109 -338
rect -159 -378 -97 -372
rect -31 -378 31 -372
rect 97 -378 159 -372
<< pwell >>
rect -359 -510 359 510
<< nmoslvt >>
rect -163 -300 -93 300
rect -35 -300 35 300
rect 93 -300 163 300
<< ndiff >>
rect -221 288 -163 300
rect -221 -288 -209 288
rect -175 -288 -163 288
rect -221 -300 -163 -288
rect -93 288 -35 300
rect -93 -288 -81 288
rect -47 -288 -35 288
rect -93 -300 -35 -288
rect 35 288 93 300
rect 35 -288 47 288
rect 81 -288 93 288
rect 35 -300 93 -288
rect 163 288 221 300
rect 163 -288 175 288
rect 209 -288 221 288
rect 163 -300 221 -288
<< ndiffc >>
rect -209 -288 -175 288
rect -81 -288 -47 288
rect 47 -288 81 288
rect 175 -288 209 288
<< psubdiff >>
rect -323 440 -227 474
rect 227 440 323 474
rect -323 378 -289 440
rect 289 378 323 440
rect -323 -440 -289 -378
rect 289 -440 323 -378
rect -323 -474 -227 -440
rect 227 -474 323 -440
<< psubdiffcont >>
rect -227 440 227 474
rect -323 -378 -289 378
rect 289 -378 323 378
rect -227 -474 227 -440
<< poly >>
rect -163 372 -93 388
rect -163 338 -147 372
rect -109 338 -93 372
rect -163 300 -93 338
rect -35 372 35 388
rect -35 338 -19 372
rect 19 338 35 372
rect -35 300 35 338
rect 93 372 163 388
rect 93 338 109 372
rect 147 338 163 372
rect 93 300 163 338
rect -163 -338 -93 -300
rect -163 -372 -147 -338
rect -109 -372 -93 -338
rect -163 -388 -93 -372
rect -35 -338 35 -300
rect -35 -372 -19 -338
rect 19 -372 35 -338
rect -35 -388 35 -372
rect 93 -338 163 -300
rect 93 -372 109 -338
rect 147 -372 163 -338
rect 93 -388 163 -372
<< polycont >>
rect -147 338 -109 372
rect -19 338 19 372
rect 109 338 147 372
rect -147 -372 -109 -338
rect -19 -372 19 -338
rect 109 -372 147 -338
<< locali >>
rect -323 440 -227 474
rect 227 440 323 474
rect -323 378 -289 440
rect 289 378 323 440
rect -163 338 -147 372
rect -109 338 -93 372
rect -35 338 -19 372
rect 19 338 35 372
rect 93 338 109 372
rect 147 338 163 372
rect -209 288 -175 304
rect -209 -304 -175 -288
rect -81 288 -47 304
rect -81 -304 -47 -288
rect 47 288 81 304
rect 47 -304 81 -288
rect 175 288 209 304
rect 175 -304 209 -288
rect -163 -372 -147 -338
rect -109 -372 -93 -338
rect -35 -372 -19 -338
rect 19 -372 35 -338
rect 93 -372 109 -338
rect 147 -372 163 -338
rect -323 -440 -289 -378
rect 289 -440 323 -378
rect -323 -474 -227 -440
rect 227 -474 323 -440
<< viali >>
rect -147 338 -109 372
rect -19 338 19 372
rect 109 338 147 372
rect -209 -288 -175 288
rect -81 -288 -47 288
rect 47 -288 81 288
rect 175 -288 209 288
rect -147 -372 -109 -338
rect -19 -372 19 -338
rect 109 -372 147 -338
<< metal1 >>
rect -159 372 -97 378
rect -159 338 -147 372
rect -109 338 -97 372
rect -159 332 -97 338
rect -31 372 31 378
rect -31 338 -19 372
rect 19 338 31 372
rect -31 332 31 338
rect 97 372 159 378
rect 97 338 109 372
rect 147 338 159 372
rect 97 332 159 338
rect -215 288 -169 300
rect -215 -288 -209 288
rect -175 -288 -169 288
rect -215 -300 -169 -288
rect -87 288 -41 300
rect -87 -288 -81 288
rect -47 -288 -41 288
rect -87 -300 -41 -288
rect 41 288 87 300
rect 41 -288 47 288
rect 81 -288 87 288
rect 41 -300 87 -288
rect 169 288 215 300
rect 169 -288 175 288
rect 209 -288 215 288
rect 169 -300 215 -288
rect -159 -338 -97 -332
rect -159 -372 -147 -338
rect -109 -372 -97 -338
rect -159 -378 -97 -372
rect -31 -338 31 -332
rect -31 -372 -19 -338
rect 19 -372 31 -338
rect -31 -378 31 -372
rect 97 -338 159 -332
rect 97 -372 109 -338
rect 147 -372 159 -338
rect 97 -378 159 -372
<< properties >>
string FIXED_BBOX -306 -457 306 457
string gencell sky130_fd_pr__nfet_01v8_lvt
string library sky130
string parameters w 3 l 0.35 m 1 nf 3 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
