magic
tech sky130A
magscale 1 2
timestamp 1666563879
<< locali >>
rect -6950 -6890 -6760 -6850
rect -6860 -6970 -6820 -6890
<< viali >>
rect -7150 -5750 -7094 -5694
rect -6650 -5750 -6594 -5694
rect -4430 -5720 -4374 -5664
rect -6870 -7700 -6814 -7644
rect -5420 -7700 -5364 -7644
rect -4700 -7700 -4644 -7644
rect -3580 -7700 -3524 -7644
<< metal1 >>
rect -3890 -3090 -3880 -3026
rect -3816 -3090 -3806 -3026
rect -6394 -3549 -6161 -3140
rect -6160 -5430 -5020 -5110
rect -7010 -5460 -5020 -5430
rect -7162 -5694 -7082 -5688
rect -6662 -5694 -6582 -5688
rect -7162 -5750 -7150 -5694
rect -7094 -5750 -7082 -5694
rect -6910 -5750 -6900 -5694
rect -6844 -5750 -6834 -5694
rect -6662 -5750 -6650 -5694
rect -6594 -5750 -6582 -5694
rect -7162 -5756 -7082 -5750
rect -6890 -5890 -6850 -5750
rect -6662 -5756 -6582 -5750
rect -7010 -5930 -6700 -5890
rect -7220 -6090 -7200 -6060
rect -7220 -6130 -7190 -6090
rect -7220 -6180 -6570 -6130
rect -7220 -6520 -7190 -6180
rect -7150 -6490 -7070 -6440
rect -6620 -6490 -6550 -6440
rect -7220 -6600 -7200 -6520
rect -6520 -6580 -6490 -6020
rect -6438 -6340 -6428 -6288
rect -7060 -6640 -6640 -6600
rect -7320 -6800 -7100 -6750
rect -6890 -7040 -6850 -6640
rect -6620 -6766 -6550 -6750
rect -6370 -6766 -6340 -5460
rect -6160 -5610 -5020 -5460
rect -4350 -5658 -4300 -3380
rect -4442 -5664 -4320 -5658
rect -4442 -5720 -4430 -5664
rect -4374 -5710 -4320 -5664
rect -4268 -5710 -4258 -5658
rect -4374 -5720 -4300 -5710
rect -4442 -5726 -4300 -5720
rect -4700 -5960 -4690 -5896
rect -4626 -5960 -4616 -5896
rect -6620 -6796 -6340 -6766
rect -6620 -6800 -6550 -6796
rect -7040 -7080 -6690 -7040
rect -7090 -7300 -7080 -7288
rect -7510 -7340 -7080 -7300
rect -7028 -7300 -7018 -7288
rect -6900 -7300 -6890 -7130
rect -6830 -7300 -6800 -7130
rect -6670 -7300 -6660 -7288
rect -7028 -7340 -6660 -7300
rect -6608 -7300 -6598 -7288
rect -6608 -7340 -6500 -7300
rect -6900 -7520 -6890 -7340
rect -6830 -7520 -6800 -7340
rect -7100 -7660 -7060 -7570
rect -6882 -7644 -6802 -7638
rect -6882 -7660 -6870 -7644
rect -7200 -7700 -6870 -7660
rect -6814 -7660 -6802 -7644
rect -6670 -7660 -6630 -7560
rect -6814 -7700 -6510 -7660
rect -6882 -7706 -6802 -7700
rect -6140 -7760 -5820 -7150
rect -4700 -7240 -4690 -7188
rect -4638 -7240 -4628 -7188
rect -4350 -7510 -4300 -5726
rect -4680 -7590 -4240 -7550
rect -4230 -7560 -4190 -3330
rect -4120 -3580 -4070 -3380
rect -3880 -3580 -3810 -3090
rect -4120 -3630 -3810 -3580
rect -4120 -3970 -4070 -3630
rect -3880 -3970 -3810 -3630
rect -4120 -4020 -3800 -3970
rect -4120 -5670 -4070 -4020
rect -3880 -5670 -3810 -4020
rect -4120 -5720 -3800 -5670
rect -4120 -6570 -4070 -5720
rect -3880 -6570 -3810 -5720
rect -4120 -6620 -3800 -6570
rect -4120 -7410 -4070 -6620
rect -3880 -7410 -3810 -6620
rect -3610 -7280 -3560 -3500
rect -3620 -7298 -3520 -7280
rect -3620 -7350 -3610 -7298
rect -3558 -7300 -3520 -7298
rect -3558 -7350 -3548 -7300
rect -4120 -7460 -3800 -7410
rect -4120 -7510 -4070 -7460
rect -3880 -7540 -3810 -7460
rect -3610 -7550 -3560 -7350
rect -3314 -7544 -3244 -3550
rect -3314 -7600 -3300 -7544
rect -3244 -7600 -3234 -7544
rect -5432 -7644 -5352 -7638
rect -5432 -7700 -5420 -7644
rect -5364 -7700 -5352 -7644
rect -5432 -7706 -5352 -7700
rect -4712 -7644 -4632 -7638
rect -4712 -7700 -4700 -7644
rect -4644 -7700 -4632 -7644
rect -4712 -7706 -4632 -7700
rect -3592 -7644 -3512 -7638
rect -3592 -7700 -3580 -7644
rect -3524 -7700 -3512 -7644
rect -3592 -7706 -3512 -7700
<< via1 >>
rect -3880 -3090 -3816 -3026
rect -7150 -5750 -7094 -5694
rect -6900 -5750 -6844 -5694
rect -6650 -5750 -6594 -5694
rect -6490 -6340 -6438 -6288
rect -4430 -5720 -4374 -5664
rect -4320 -5710 -4268 -5658
rect -4690 -5960 -4626 -5896
rect -7080 -7340 -7028 -7288
rect -6660 -7340 -6608 -7288
rect -6870 -7700 -6814 -7644
rect -4690 -7240 -4638 -7188
rect -3610 -7350 -3558 -7298
rect -3300 -7600 -3244 -7544
rect -5420 -7700 -5364 -7644
rect -4700 -7700 -4644 -7644
rect -3580 -7700 -3524 -7644
<< metal2 >>
rect -3880 -3026 -3816 -3016
rect -3880 -3100 -3816 -3090
rect -4320 -5650 -4268 -5648
rect -7320 -5658 -3970 -5650
rect -7320 -5664 -4320 -5658
rect -7320 -5694 -4430 -5664
rect -7320 -5750 -7150 -5694
rect -7094 -5750 -6900 -5694
rect -6844 -5750 -6650 -5694
rect -6594 -5720 -4430 -5694
rect -4374 -5710 -4320 -5664
rect -4268 -5710 -3970 -5658
rect -4374 -5720 -3970 -5710
rect -6594 -5750 -3970 -5720
rect -7320 -5770 -3970 -5750
rect -4690 -5896 -4626 -5886
rect -4690 -5970 -4626 -5960
rect -6490 -6288 -6438 -6278
rect -6438 -6340 -4820 -6290
rect -6490 -6350 -6438 -6340
rect -4870 -7190 -4820 -6340
rect -4690 -7188 -4638 -7178
rect -4870 -7240 -4690 -7190
rect -4690 -7250 -4638 -7240
rect -7080 -7288 -7028 -7278
rect -7100 -7340 -7080 -7300
rect -6660 -7288 -6608 -7278
rect -7028 -7340 -6660 -7300
rect -3610 -7298 -3558 -7288
rect -6608 -7340 -3610 -7300
rect -7080 -7350 -7028 -7340
rect -6660 -7350 -6608 -7340
rect -3558 -7340 -3550 -7300
rect -3610 -7360 -3558 -7350
rect -3300 -7544 -3244 -7534
rect -3300 -7610 -3244 -7600
rect -6870 -7644 -6814 -7634
rect -6870 -7710 -6814 -7700
rect -5420 -7644 -5364 -7634
rect -5420 -7710 -5364 -7700
rect -4700 -7644 -4644 -7634
rect -4700 -7710 -4644 -7700
rect -3580 -7644 -3524 -7634
rect -3580 -7710 -3524 -7700
<< via2 >>
rect -3880 -3090 -3816 -3026
rect -4690 -5960 -4626 -5896
rect -3300 -7600 -3244 -7544
rect -6870 -7700 -6814 -7644
rect -5420 -7700 -5364 -7644
rect -4700 -7700 -4644 -7644
rect -3580 -7700 -3524 -7644
<< metal3 >>
rect -8020 -2160 -2721 17840
rect -3900 -3026 -3750 -3020
rect -3900 -3090 -3880 -3026
rect -3816 -3090 -3750 -3026
rect -3900 -3100 -3750 -3090
rect -4700 -5896 -4610 -5830
rect -4700 -5960 -4690 -5896
rect -4626 -5960 -4610 -5896
rect -4700 -5970 -4610 -5960
rect -3310 -7544 -3234 -7539
rect -3310 -7600 -3300 -7544
rect -3244 -7600 -3234 -7544
rect -7340 -7644 -3170 -7600
rect -7340 -7700 -6870 -7644
rect -6814 -7700 -5420 -7644
rect -5364 -7700 -4700 -7644
rect -4644 -7700 -3580 -7644
rect -3524 -7700 -3170 -7644
rect -7340 -7740 -3170 -7700
<< via3 >>
rect -3880 -3090 -3816 -3026
rect -4690 -5960 -4626 -5896
<< metal4 >>
rect -5550 -2960 -4610 -2870
rect -4700 -5896 -4610 -2960
rect -2848 -3020 -2748 -2960
rect -3900 -3026 -2748 -3020
rect -3900 -3090 -3880 -3026
rect -3816 -3090 -2748 -3026
rect -3900 -3100 -2748 -3090
rect -4700 -5960 -4690 -5896
rect -4626 -5960 -4610 -5896
rect -4700 -5970 -4610 -5960
use sky130_fd_pr__cap_mim_m3_1_L4YDVW  XC4
timestamp 1662478139
transform 1 0 -5370 0 1 7640
box -2650 -10600 2649 10600
use sky130_fd_pr__nfet_01v8_lvt_EA9ZG2  XM54
timestamp 1662478139
transform 1 0 -7131 0 1 -6620
box -221 -310 221 310
use sky130_fd_pr__nfet_01v8_lvt_EA9ZG2  XM55
timestamp 1662478139
transform 1 0 -6579 0 1 -6620
box -221 -310 221 310
use sky130_fd_pr__nfet_01v8_lvt_BSMWRE  XM56
timestamp 1662478139
transform 0 1 -6853 -1 0 -7326
box -396 -519 396 519
use sky130_fd_pr__nfet_01v8_lvt_F8HAAN  XM57
timestamp 1662478139
transform 1 0 -3566 0 1 -5531
box -396 -2191 396 2191
use sky130_fd_pr__pfet_01v8_lvt_X3YSY6  XM58
timestamp 1662478139
transform 1 0 -6612 0 1 -5991
box -246 -319 246 319
use sky130_fd_pr__pfet_01v8_lvt_X3YSY6  XM59
timestamp 1662478139
transform 1 0 -7104 0 1 -5991
box -246 -319 246 319
use sky130_fd_pr__pfet_01v8_lvt_ER7KZU  XM60
timestamp 1662478139
transform 1 0 -4208 0 1 -5441
box -246 -2281 246 2281
use sky130_fd_pr__res_high_po_0p35_ZMQPMJ  XR34
timestamp 1662478139
transform 1 0 -4655 0 1 -6724
box -201 -998 201 998
use sky130_fd_pr__res_xhigh_po_5p73_Q3K92U  XR35
timestamp 1662478139
transform 1 0 -5595 0 1 -6532
box -739 -1190 739 1190
use sky130_fd_pr__res_xhigh_po_5p73_Q3K92U  XR37
timestamp 1662478139
transform 1 0 -5595 0 1 -4152
box -739 -1190 739 1190
<< labels >>
rlabel metal2 -7300 -5650 -7300 -5650 1 vdd
port 6 n
rlabel metal3 -7188 -7740 -7188 -7740 5 vss
port 5 s
rlabel metal1 -6020 -7760 -6020 -7760 5 vinn
port 1 s
rlabel metal1 -7320 -6770 -7320 -6770 7 vref
port 2 w
rlabel metal1 -7510 -7320 -7510 -7320 7 vbcm
port 4 w
rlabel metal1 -6394 -3420 -6394 -3420 7 vinp
port 0 w
rlabel metal1 -7010 -5440 -7010 -5440 7 vcm
rlabel metal4 -2748 -3070 -2748 -3070 1 vc
port 3 n
<< end >>
