magic
tech sky130A
magscale 1 2
timestamp 1672090405
<< locali >>
rect 12696 -754 12730 -612
rect 16764 -754 16798 -612
rect 14870 -1372 14906 -1234
rect 9156 -1586 9702 -1550
rect 19044 -1660 19724 -1622
rect 14766 -1838 14904 -1802
rect 10280 -1886 11422 -1850
rect 11998 -1888 12642 -1850
rect 17018 -1886 17252 -1852
rect 17828 -1886 18468 -1848
rect 12718 -2400 12752 -2260
rect 13500 -2400 13534 -2260
rect 13804 -2400 13838 -2260
rect 14992 -2400 15324 -2366
rect 15610 -2400 16124 -2366
rect 13176 -2770 13232 -2758
rect 13176 -2898 13184 -2770
rect 13224 -2898 13232 -2770
rect 13176 -2902 13232 -2898
rect 15598 -2776 15654 -2770
rect 15598 -2906 15604 -2776
rect 15650 -2906 15654 -2776
rect 15598 -2914 15654 -2906
<< viali >>
rect 13184 -2898 13224 -2770
rect 15604 -2906 15650 -2776
<< metal1 >>
rect 8980 -550 12076 -504
rect 14660 -550 19904 -504
rect 8980 -1178 9046 -550
rect 10102 -1172 18646 -1124
rect 10102 -1480 10168 -1172
rect 11824 -1480 17428 -1432
rect 12540 -2200 16302 -2152
rect 12540 -2508 12606 -2200
rect 13166 -2768 13232 -2758
rect 13166 -2906 13176 -2768
rect 13228 -2906 13232 -2768
rect 15590 -2772 15662 -2762
rect 13326 -2812 15502 -2778
rect 13166 -2916 13232 -2906
rect 15132 -4042 15172 -2812
rect 15590 -2906 15596 -2772
rect 15654 -2906 15662 -2772
rect 15590 -2918 15662 -2906
rect 15796 -4048 15834 -2200
rect 16236 -2502 16302 -2200
rect 17112 -4036 17154 -1480
rect 18104 -4056 18142 -1172
rect 18580 -1472 18646 -1172
rect 19342 -4040 19380 -550
rect 19838 -1258 19904 -550
<< via1 >>
rect 13176 -2770 13228 -2768
rect 13176 -2898 13184 -2770
rect 13184 -2898 13224 -2770
rect 13224 -2898 13228 -2770
rect 13176 -2906 13228 -2898
rect 15596 -2776 15654 -2772
rect 15596 -2906 15604 -2776
rect 15604 -2906 15650 -2776
rect 15650 -2906 15654 -2776
<< metal2 >>
rect 9374 -1338 11938 -1330
rect 8452 -1350 11938 -1338
rect 8452 -1520 11720 -1350
rect 11902 -1520 11938 -1350
rect 17314 -1346 19522 -1330
rect 8452 -1578 11938 -1520
rect 17314 -1522 17608 -1346
rect 17844 -1418 19522 -1346
rect 17844 -1522 20432 -1418
rect 17314 -1578 20432 -1522
rect 8452 -1586 9578 -1578
rect 19326 -1666 20432 -1578
rect 13146 -2668 13280 -2538
rect 15542 -2668 15680 -2538
rect 12470 -2768 13306 -2668
rect 12470 -2906 13176 -2768
rect 13228 -2906 13306 -2768
rect 12470 -2916 13306 -2906
rect 15542 -2772 16378 -2668
rect 15542 -2906 15596 -2772
rect 15654 -2906 16378 -2772
rect 15542 -2916 16378 -2906
<< via2 >>
rect 12002 -324 12232 -198
rect 17562 -544 17800 -426
rect 8468 -1256 8688 -1134
rect 11720 -1520 11902 -1350
rect 20204 -1338 20416 -1234
rect 16704 -1564 16928 -1456
rect 17608 -1522 17844 -1346
rect 9978 -1770 10186 -1658
rect 11726 -1758 11912 -1672
rect 14990 -1762 15214 -1654
rect 17334 -1744 17474 -1682
rect 18556 -1762 18760 -1664
rect 12742 -1970 12960 -1874
rect 14442 -2176 14678 -2062
<< metal3 >>
rect 8452 -198 12248 -184
rect 8452 -324 12002 -198
rect 12232 -324 12248 -198
rect 8452 -338 12248 -324
rect 8452 -1122 8606 -338
rect 17542 -426 20426 -408
rect 17542 -544 17562 -426
rect 17800 -544 20426 -426
rect 17542 -560 20426 -544
rect 10024 -956 13052 -804
rect 8452 -1134 8702 -1122
rect 8452 -1136 8468 -1134
rect 8452 -1264 8462 -1136
rect 8688 -1256 8702 -1134
rect 8596 -1264 8702 -1256
rect 8452 -1274 8702 -1264
rect 8452 -1276 8606 -1274
rect 10024 -1646 10216 -956
rect 16442 -1180 18722 -1028
rect 11692 -1350 11936 -1328
rect 11692 -1520 11720 -1350
rect 11902 -1520 11936 -1350
rect 17580 -1346 17862 -1328
rect 11692 -1542 11936 -1520
rect 16678 -1456 17496 -1442
rect 16678 -1564 16704 -1456
rect 16928 -1564 17496 -1456
rect 17580 -1522 17608 -1346
rect 17844 -1522 17862 -1346
rect 17580 -1542 17862 -1522
rect 16678 -1584 17496 -1564
rect 9962 -1658 10216 -1646
rect 9962 -1770 9978 -1658
rect 10208 -1768 10216 -1658
rect 10186 -1770 10216 -1768
rect 9962 -1784 10216 -1770
rect 11538 -1652 15232 -1640
rect 11538 -1768 11554 -1652
rect 11722 -1654 15232 -1652
rect 11722 -1672 14990 -1654
rect 11722 -1758 11726 -1672
rect 11912 -1758 14990 -1672
rect 11722 -1762 14990 -1758
rect 15214 -1762 15232 -1654
rect 11722 -1768 15232 -1762
rect 11538 -1780 15232 -1768
rect 17314 -1660 17496 -1584
rect 17314 -1758 17328 -1660
rect 17484 -1758 17496 -1660
rect 17314 -1778 17496 -1758
rect 18532 -1644 18722 -1180
rect 20274 -1210 20426 -560
rect 20174 -1224 20426 -1210
rect 20174 -1234 20288 -1224
rect 20412 -1234 20426 -1224
rect 20174 -1338 20204 -1234
rect 20416 -1338 20426 -1234
rect 20174 -1346 20288 -1338
rect 20412 -1346 20426 -1338
rect 20174 -1362 20426 -1346
rect 18532 -1656 18844 -1644
rect 18532 -1664 18664 -1656
rect 18532 -1762 18556 -1664
rect 18532 -1784 18664 -1762
rect 18828 -1784 18844 -1656
rect 18532 -1796 18844 -1784
rect 5100 -2240 7800 -1840
rect 12714 -1874 12990 -1850
rect 12714 -1970 12742 -1874
rect 12960 -1970 12990 -1874
rect 12714 -1990 12990 -1970
rect 5100 -3040 12000 -2240
rect 12776 -2476 12990 -1990
rect 14424 -2062 16108 -2048
rect 14424 -2176 14442 -2062
rect 14678 -2176 16108 -2062
rect 14424 -2188 16108 -2176
rect 12394 -2486 12990 -2476
rect 12394 -2598 12800 -2486
rect 12980 -2598 12990 -2486
rect 14648 -2468 15440 -2450
rect 12394 -2612 12990 -2598
rect 12776 -2614 12990 -2612
rect 13120 -2556 13334 -2540
rect 13120 -2724 13138 -2556
rect 13306 -2724 13334 -2556
rect 14648 -2566 14780 -2468
rect 14932 -2566 15440 -2468
rect 15894 -2472 16108 -2188
rect 15894 -2486 16446 -2472
rect 14648 -2610 15440 -2566
rect 15536 -2554 15750 -2538
rect 13120 -2740 13334 -2724
rect 13400 -2698 14178 -2670
rect 13400 -2802 13916 -2698
rect 14090 -2802 14178 -2698
rect 15536 -2728 15546 -2554
rect 15736 -2728 15750 -2554
rect 15894 -2596 15916 -2486
rect 16094 -2596 16446 -2486
rect 15894 -2612 16446 -2596
rect 15536 -2740 15750 -2728
rect 13400 -2830 14178 -2802
rect 16968 -3040 19667 -2240
rect 20980 -3040 21210 -2240
rect 5100 -4040 14218 -3040
rect 14518 -4040 23779 -3040
<< via3 >>
rect 8462 -1256 8468 -1136
rect 8468 -1256 8596 -1136
rect 8462 -1264 8596 -1256
rect 11720 -1520 11902 -1350
rect 17608 -1522 17844 -1346
rect 10040 -1768 10186 -1658
rect 10186 -1768 10208 -1658
rect 11554 -1768 11722 -1652
rect 17328 -1682 17484 -1660
rect 17328 -1744 17334 -1682
rect 17334 -1744 17474 -1682
rect 17474 -1744 17484 -1682
rect 17328 -1758 17484 -1744
rect 20288 -1234 20412 -1224
rect 20288 -1338 20412 -1234
rect 20288 -1346 20412 -1338
rect 18664 -1664 18828 -1656
rect 18664 -1762 18760 -1664
rect 18760 -1762 18828 -1664
rect 18664 -1784 18828 -1762
rect 12800 -2598 12980 -2486
rect 13138 -2724 13306 -2556
rect 14780 -2566 14932 -2468
rect 13916 -2802 14090 -2698
rect 15546 -2728 15736 -2554
rect 15916 -2596 16094 -2486
<< metal4 >>
rect 7466 -1136 8606 -1122
rect 7466 -1264 8462 -1136
rect 8596 -1264 8606 -1136
rect 7466 -1276 8606 -1264
rect 20274 -1224 21956 -1210
rect 11692 -1346 17862 -1328
rect 11692 -1350 17608 -1346
rect 11692 -1520 11720 -1350
rect 11902 -1520 17608 -1350
rect 11692 -1522 17608 -1520
rect 17844 -1522 17862 -1346
rect 20274 -1346 20288 -1224
rect 20412 -1346 21956 -1224
rect 20274 -1362 21956 -1346
rect 11692 -1542 17862 -1522
rect 10024 -1658 10216 -1646
rect 10024 -1768 10040 -1658
rect 10208 -1768 10216 -1658
rect 10024 -2514 10216 -1768
rect 11538 -1652 11732 -1640
rect 11538 -1768 11554 -1652
rect 11722 -1768 11732 -1652
rect 11538 -2470 11732 -1768
rect 12776 -2486 12990 -2474
rect 12776 -2598 12800 -2486
rect 12980 -2598 12990 -2486
rect 12776 -3268 12990 -2598
rect 13120 -2556 13334 -1542
rect 13120 -2724 13138 -2556
rect 13306 -2724 13334 -2556
rect 14740 -2468 14964 -2450
rect 14740 -2566 14780 -2468
rect 14932 -2566 14964 -2468
rect 13120 -2740 13334 -2724
rect 13896 -2698 14110 -2676
rect 13896 -2802 13916 -2698
rect 14090 -2802 14110 -2698
rect 13896 -3324 14110 -2802
rect 14740 -3258 14964 -2566
rect 15536 -2554 15750 -1542
rect 17304 -1660 17496 -1646
rect 17304 -1758 17328 -1660
rect 17484 -1758 17496 -1660
rect 17304 -2420 17496 -1758
rect 18650 -1656 18844 -1644
rect 18650 -1784 18664 -1656
rect 18828 -1784 18844 -1656
rect 18650 -2466 18844 -1784
rect 15536 -2728 15546 -2554
rect 15736 -2728 15750 -2554
rect 15536 -2740 15750 -2728
rect 15894 -2486 16108 -2472
rect 15894 -2596 15916 -2486
rect 16094 -2596 16108 -2486
rect 15894 -3244 16108 -2596
use sky130_fd_pr__cap_mim_m3_1_3ZFDVT  XC1 /foss/designs/layout
timestamp 1671746299
transform -1 0 13827 0 1 -3540
box -450 -500 449 500
use sky130_fd_pr__cap_mim_m3_1_VCH7EQ  XC2 /foss/designs/layout
timestamp 1671746277
transform -1 0 12627 0 1 -3540
box -750 -500 749 500
use sky130_fd_pr__cap_mim_m3_1_MYMY8D  XC3 /foss/designs/layout
timestamp 1671746242
transform -1 0 11127 0 1 -3140
box -750 -900 749 900
use sky130_fd_pr__cap_mim_m3_1_CYFFME  XC4 /foss/designs/layout
timestamp 1671746218
transform -1 0 9027 0 1 -3140
box -1350 -900 1349 900
use sky130_fd_pr__cap_mim_m3_1_A6B8BZ  XC5 /foss/designs/layout
timestamp 1671746188
transform -1 0 6327 0 1 -2340
box -1350 -1700 1349 1700
use sky130_fd_pr__cap_mim_m3_1_3ZFDVT  XC6
timestamp 1671746299
transform 1 0 15052 0 1 -3540
box -450 -500 449 500
use sky130_fd_pr__cap_mim_m3_1_VCH7EQ  XC7
timestamp 1671746277
transform 1 0 16254 0 1 -3540
box -750 -500 749 500
use sky130_fd_pr__cap_mim_m3_1_MYMY8D  XC8
timestamp 1671746242
transform 1 0 17754 0 1 -3140
box -750 -900 749 900
use sky130_fd_pr__cap_mim_m3_1_CYFFME  XC9
timestamp 1671746218
transform 1 0 19854 0 1 -3140
box -1350 -900 1349 900
use sky130_fd_pr__cap_mim_m3_1_A6B8BZ  XC10
timestamp 1671746188
transform 1 0 22554 0 1 -2340
box -1350 -1700 1349 1700
use sky130_fd_pr__nfet_01v8_lvt_648S5X  XM1 /foss/designs/layout
timestamp 1671770132
transform 1 0 13360 0 1 -2640
box -212 -310 210 310
use sky130_fd_pr__nfet_01v8_lvt_DJ7QE5  XM2 /foss/designs/layout
timestamp 1671754502
transform 1 0 12526 0 1 -2640
box -264 -310 262 310
use sky130_fd_pr__nfet_01v8_lvt_HNLS5R  XM3 /foss/designs/layout
timestamp 1671762831
transform 1 0 11714 0 1 -1612
box -360 -310 358 310
use sky130_fd_pr__nfet_01v8_lvt_HNLS5R  XM4
timestamp 1671762831
transform 1 0 9992 0 1 -1612
box -360 -310 358 310
use sky130_fd_pr__nfet_01v8_lvt_B6HS5D  XM5 /foss/designs/layout
timestamp 1671768516
transform 1 0 8774 0 1 -1310
box -456 -310 454 310
use sky130_fd_pr__nfet_01v8_lvt_648S5X  XM6
timestamp 1671770132
transform -1 0 15468 0 1 -2640
box -212 -310 210 310
use sky130_fd_pr__nfet_01v8_lvt_DJ7QE5  XM7
timestamp 1671754502
transform -1 0 16316 0 1 -2640
box -264 -310 262 310
use sky130_fd_pr__nfet_01v8_lvt_HNLS5R  XM8
timestamp 1671762831
transform -1 0 17538 0 1 -1612
box -360 -310 358 310
use sky130_fd_pr__nfet_01v8_lvt_HNLS5R  XM9
timestamp 1671762831
transform -1 0 18756 0 1 -1610
box -360 -310 358 310
use sky130_fd_pr__nfet_01v8_lvt_B6HS5D  XM10
timestamp 1671768516
transform -1 0 20110 0 1 -1390
box -456 -310 454 310
use sky130_fd_pr__nfet_01v8_lvt_9DHFGX  XM11 /foss/designs/layout
timestamp 1671754915
transform 1 0 14417 0 1 -2640
box -648 -310 647 310
use sky130_fd_pr__nfet_01v8_lvt_YTLFGX  XM12 /foss/designs/layout
timestamp 1671827388
transform 1 0 13708 0 1 -2020
box -1128 -310 1126 310
use sky130_fd_pr__nfet_01v8_lvt_YTLFGX  XM13
timestamp 1671827388
transform 1 0 15962 0 -1 -1612
box -1128 -310 1126 310
use sky130_fd_pr__nfet_01v8_lvt_A33GGX  XM14 /foss/designs/layout
timestamp 1671764736
transform 1 0 14748 0 1 -992
box -2088 -310 2086 310
use sky130_fd_pr__nfet_01v8_lvt_LELFGX  XM15 /foss/designs/layout
timestamp 1671767400
transform 1 0 14902 0 1 -372
box -3048 -310 3046 310
<< labels >>
flabel metal4 11902 -1542 17608 -1328 0 FreeSans 800 0 0 0 GND
flabel metal1 15132 -4042 15172 -2778 0 FreeSans 800 0 0 0 ctrll1
flabel metal1 15796 -4048 15834 -2152 0 FreeSans 800 0 0 0 ctrll2
flabel metal1 17112 -4036 17154 -1432 0 FreeSans 800 0 0 0 ctrll3
flabel metal1 18104 -4056 18142 -1124 0 FreeSans 800 0 0 0 ctrll4
flabel metal1 19342 -4040 19380 -504 0 FreeSans 800 0 0 0 ctrll5
flabel space 5100 -4040 14399 -3040 0 FreeSans 800 0 0 0 IN2
flabel space 14480 -4040 23779 -3040 0 FreeSans 800 0 0 0 IN
<< end >>
