magic
tech sky130A
magscale 1 2
timestamp 1672483164
<< pwell >>
rect 53403 -7310 53408 -7308
<< ndiff >>
rect 53403 -7310 53408 -7308
<< locali >>
rect 64128 -5922 64180 -5920
rect 51840 -5960 64180 -5922
rect 51840 -6120 51896 -5960
rect 52286 -6008 52336 -5960
rect 52668 -6010 52718 -5960
rect 53050 -6010 53100 -5960
rect 53434 -6010 53484 -5960
rect 53818 -6006 53868 -5960
rect 54204 -6008 54254 -5960
rect 54584 -6010 54634 -5960
rect 54970 -6010 55020 -5960
rect 55356 -6008 55406 -5960
rect 55736 -6010 55786 -5960
rect 56120 -6012 56170 -5960
rect 56508 -6010 56558 -5960
rect 56888 -6010 56938 -5960
rect 57272 -6010 57322 -5960
rect 57658 -6010 57708 -5960
rect 58474 -6008 58524 -5960
rect 58860 -6010 58910 -5960
rect 59246 -6012 59296 -5960
rect 59630 -6010 59680 -5960
rect 60012 -6012 60062 -5960
rect 60398 -6010 60448 -5960
rect 60782 -6008 60832 -5960
rect 61164 -6008 61214 -5960
rect 61550 -6010 61600 -5960
rect 61932 -6008 61982 -5960
rect 62316 -6010 62366 -5960
rect 62698 -6010 62748 -5960
rect 63084 -6010 63134 -5960
rect 63466 -6008 63516 -5960
rect 63852 -6006 63902 -5960
rect 51840 -6176 51842 -6120
rect 64128 -6176 64180 -5960
rect 51840 -6372 51896 -6176
rect 51998 -6372 52042 -6306
rect 52380 -6372 52424 -6306
rect 52766 -6372 52810 -6304
rect 53154 -6372 53198 -6312
rect 53536 -6372 53580 -6312
rect 53916 -6372 53960 -6314
rect 54304 -6372 54348 -6310
rect 54688 -6372 54732 -6310
rect 55078 -6372 55122 -6304
rect 55454 -6372 55498 -6310
rect 55840 -6372 55884 -6310
rect 56218 -6372 56262 -6314
rect 56606 -6372 56650 -6308
rect 56988 -6372 57032 -6314
rect 57382 -6372 57426 -6312
rect 57756 -6372 57800 -6308
rect 58188 -6372 58232 -6308
rect 58574 -6372 58618 -6308
rect 58962 -6372 59006 -6314
rect 59344 -6372 59388 -6318
rect 59726 -6372 59770 -6314
rect 60112 -6372 60156 -6310
rect 60492 -6372 60536 -6314
rect 60878 -6372 60922 -6318
rect 61266 -6372 61310 -6316
rect 61654 -6372 61698 -6308
rect 62034 -6372 62078 -6314
rect 62418 -6372 62462 -6314
rect 62796 -6372 62840 -6312
rect 63182 -6372 63226 -6312
rect 63566 -6372 63610 -6314
rect 63958 -6372 64002 -6316
rect 64128 -6372 64180 -6232
rect 48302 -6542 48426 -6396
rect 51840 -6408 64180 -6372
rect 51858 -6410 64180 -6408
rect 51732 -6534 64248 -6500
rect 51732 -7036 51772 -6534
rect 52292 -6624 52336 -6534
rect 52666 -6624 52710 -6534
rect 53056 -6624 53100 -6534
rect 53438 -6624 53482 -6534
rect 53822 -6624 53866 -6534
rect 54212 -6620 54256 -6534
rect 54584 -6624 54628 -6534
rect 54970 -6624 55014 -6534
rect 55360 -6630 55404 -6534
rect 55740 -6626 55784 -6534
rect 56122 -6626 56166 -6534
rect 56502 -6622 56546 -6534
rect 56890 -6620 56934 -6534
rect 57270 -6618 57314 -6534
rect 57654 -6626 57698 -6534
rect 58460 -6616 58504 -6534
rect 58844 -6616 58888 -6534
rect 59228 -6622 59272 -6534
rect 59612 -6612 59656 -6534
rect 59994 -6614 60038 -6534
rect 60386 -6620 60430 -6534
rect 60770 -6616 60814 -6534
rect 61148 -6618 61192 -6534
rect 61534 -6616 61578 -6534
rect 61922 -6622 61966 -6534
rect 62300 -6620 62344 -6534
rect 62686 -6620 62730 -6534
rect 63072 -6616 63116 -6534
rect 63460 -6620 63504 -6534
rect 63850 -6622 63894 -6534
rect 52188 -7036 52250 -6936
rect 52580 -7036 52636 -6942
rect 52962 -7036 53018 -6940
rect 53344 -7036 53400 -6942
rect 53734 -7036 53790 -6940
rect 54118 -7036 54174 -6940
rect 54498 -7036 54554 -6932
rect 54884 -7036 54940 -6944
rect 55270 -7036 55326 -6942
rect 55646 -7036 55702 -6948
rect 56030 -7036 56086 -6946
rect 56420 -7036 56476 -6948
rect 56798 -7036 56854 -6940
rect 57188 -7036 57244 -6946
rect 57566 -7036 57622 -6944
rect 58368 -7036 58424 -6942
rect 58762 -7036 58818 -6942
rect 59148 -6948 59204 -6942
rect 59138 -7036 59204 -6948
rect 59528 -7036 59584 -6940
rect 59912 -7036 59968 -6938
rect 60290 -7036 60346 -6940
rect 60676 -7036 60732 -6938
rect 61064 -7036 61120 -6942
rect 61438 -7036 61494 -6938
rect 61824 -7036 61880 -6938
rect 62218 -7036 62274 -6936
rect 62588 -7036 62644 -6940
rect 62974 -7036 63030 -6938
rect 63368 -7036 63424 -6942
rect 63742 -7036 63798 -6938
rect 64208 -7036 64248 -6534
rect 68132 -6542 68246 -6400
rect 51732 -7070 64248 -7036
<< viali >>
rect 48286 -5236 48458 -5178
rect 49920 -5280 66568 -5188
rect 68070 -5236 68242 -5178
rect 51842 -6176 51898 -6120
rect 64128 -6232 64184 -6176
rect 48274 -7764 48446 -7706
rect 49940 -7756 66588 -7664
rect 68120 -7768 68292 -7710
<< metal1 >>
rect 48274 -5178 48470 -5172
rect 47250 -6264 47260 -5190
rect 47620 -6264 47630 -5190
rect 48274 -5236 48286 -5178
rect 48458 -5236 48470 -5178
rect 68058 -5178 68254 -5172
rect 48274 -5242 48470 -5236
rect 49908 -5188 66580 -5182
rect 49908 -5280 49920 -5188
rect 66568 -5280 66580 -5188
rect 68058 -5236 68070 -5178
rect 68242 -5236 68254 -5178
rect 68058 -5242 68254 -5236
rect 49908 -5286 66580 -5280
rect 48190 -5686 48550 -5300
rect 48188 -6296 48550 -5686
rect 49880 -5400 66630 -5370
rect 49880 -5680 49910 -5400
rect 50077 -5494 50087 -5442
rect 50139 -5494 50149 -5442
rect 50267 -5493 50277 -5441
rect 50329 -5493 50339 -5441
rect 50460 -5496 50470 -5444
rect 50522 -5496 50532 -5444
rect 50652 -5491 50662 -5439
rect 50714 -5491 50724 -5439
rect 50844 -5495 50854 -5443
rect 50906 -5495 50916 -5443
rect 51036 -5490 51046 -5438
rect 51098 -5490 51108 -5438
rect 51228 -5491 51238 -5439
rect 51290 -5491 51300 -5439
rect 51418 -5490 51428 -5438
rect 51480 -5490 51490 -5438
rect 51612 -5501 51622 -5449
rect 51674 -5501 51684 -5449
rect 51801 -5499 51811 -5447
rect 51863 -5499 51873 -5447
rect 51991 -5499 52001 -5447
rect 52053 -5499 52063 -5447
rect 52190 -5500 52200 -5448
rect 52252 -5500 52262 -5448
rect 52382 -5499 52392 -5447
rect 52444 -5499 52454 -5447
rect 52572 -5500 52582 -5448
rect 52634 -5500 52644 -5448
rect 52764 -5493 52774 -5441
rect 52826 -5493 52836 -5441
rect 52956 -5495 52966 -5443
rect 53018 -5495 53028 -5443
rect 53149 -5494 53159 -5442
rect 53211 -5494 53221 -5442
rect 53341 -5492 53351 -5440
rect 53403 -5492 53413 -5440
rect 53532 -5492 53542 -5440
rect 53594 -5492 53604 -5440
rect 53726 -5497 53736 -5445
rect 53788 -5497 53798 -5445
rect 53917 -5493 53927 -5441
rect 53979 -5493 53989 -5441
rect 54109 -5489 54119 -5437
rect 54171 -5489 54181 -5437
rect 54302 -5493 54312 -5441
rect 54364 -5493 54374 -5441
rect 54494 -5493 54504 -5441
rect 54556 -5493 54566 -5441
rect 54687 -5494 54697 -5442
rect 54749 -5494 54759 -5442
rect 54879 -5492 54889 -5440
rect 54941 -5492 54951 -5440
rect 55070 -5491 55080 -5439
rect 55132 -5491 55142 -5439
rect 55261 -5490 55271 -5438
rect 55323 -5490 55333 -5438
rect 55454 -5490 55464 -5438
rect 55516 -5490 55526 -5438
rect 55645 -5499 55655 -5447
rect 55707 -5499 55717 -5447
rect 55836 -5500 55846 -5448
rect 55898 -5500 55908 -5448
rect 56026 -5501 56036 -5449
rect 56088 -5501 56098 -5449
rect 56220 -5505 56230 -5453
rect 56282 -5505 56292 -5453
rect 56412 -5507 56422 -5455
rect 56474 -5507 56484 -5455
rect 56606 -5506 56616 -5454
rect 56668 -5506 56678 -5454
rect 56798 -5503 56808 -5451
rect 56860 -5503 56870 -5451
rect 56987 -5500 56997 -5448
rect 57049 -5500 57059 -5448
rect 57181 -5498 57191 -5446
rect 57243 -5498 57253 -5446
rect 57374 -5499 57384 -5447
rect 57436 -5499 57446 -5447
rect 57567 -5500 57577 -5448
rect 57629 -5500 57639 -5448
rect 57756 -5500 57766 -5448
rect 57818 -5500 57828 -5448
rect 57949 -5500 57959 -5448
rect 58011 -5500 58021 -5448
rect 58141 -5500 58151 -5448
rect 58203 -5500 58213 -5448
rect 58332 -5500 58342 -5448
rect 58394 -5500 58404 -5448
rect 58525 -5500 58535 -5448
rect 58587 -5500 58597 -5448
rect 58716 -5499 58726 -5447
rect 58778 -5499 58788 -5447
rect 58911 -5500 58921 -5448
rect 58973 -5500 58983 -5448
rect 59100 -5500 59110 -5448
rect 59162 -5500 59172 -5448
rect 59293 -5500 59303 -5448
rect 59355 -5500 59365 -5448
rect 59485 -5500 59495 -5448
rect 59547 -5500 59557 -5448
rect 59676 -5500 59686 -5448
rect 59738 -5500 59748 -5448
rect 59868 -5500 59878 -5448
rect 59930 -5500 59940 -5448
rect 60061 -5500 60071 -5448
rect 60123 -5500 60133 -5448
rect 60250 -5501 60260 -5449
rect 60312 -5501 60322 -5449
rect 60444 -5500 60454 -5448
rect 60506 -5500 60516 -5448
rect 60635 -5500 60645 -5448
rect 60697 -5500 60707 -5448
rect 60828 -5500 60838 -5448
rect 60890 -5500 60900 -5448
rect 61020 -5500 61030 -5448
rect 61082 -5500 61092 -5448
rect 61212 -5501 61222 -5449
rect 61274 -5501 61284 -5449
rect 61405 -5499 61415 -5447
rect 61467 -5499 61477 -5447
rect 61595 -5499 61605 -5447
rect 61657 -5499 61667 -5447
rect 61788 -5501 61798 -5449
rect 61850 -5501 61860 -5449
rect 61980 -5500 61990 -5448
rect 62042 -5500 62052 -5448
rect 62173 -5499 62183 -5447
rect 62235 -5499 62245 -5447
rect 62364 -5499 62374 -5447
rect 62426 -5499 62436 -5447
rect 62556 -5500 62566 -5448
rect 62618 -5500 62628 -5448
rect 62747 -5500 62757 -5448
rect 62809 -5500 62819 -5448
rect 62939 -5500 62949 -5448
rect 63001 -5500 63011 -5448
rect 63133 -5499 63143 -5447
rect 63195 -5499 63205 -5447
rect 63325 -5500 63335 -5448
rect 63387 -5500 63397 -5448
rect 63515 -5501 63525 -5449
rect 63577 -5501 63587 -5449
rect 63706 -5502 63716 -5450
rect 63768 -5502 63778 -5450
rect 63899 -5500 63909 -5448
rect 63961 -5500 63971 -5448
rect 64092 -5499 64102 -5447
rect 64154 -5499 64164 -5447
rect 64285 -5500 64295 -5448
rect 64347 -5500 64357 -5448
rect 64476 -5500 64486 -5448
rect 64538 -5500 64548 -5448
rect 64667 -5500 64677 -5448
rect 64729 -5500 64739 -5448
rect 64860 -5500 64870 -5448
rect 64922 -5500 64932 -5448
rect 65053 -5500 65063 -5448
rect 65115 -5500 65125 -5448
rect 65244 -5500 65254 -5448
rect 65306 -5500 65316 -5448
rect 65435 -5499 65445 -5447
rect 65497 -5499 65507 -5447
rect 65626 -5499 65636 -5447
rect 65688 -5499 65698 -5447
rect 65819 -5500 65829 -5448
rect 65881 -5500 65891 -5448
rect 66013 -5500 66023 -5448
rect 66075 -5500 66085 -5448
rect 66201 -5501 66211 -5449
rect 66263 -5501 66273 -5449
rect 66395 -5509 66405 -5457
rect 66457 -5509 66467 -5457
rect 49981 -5637 49991 -5585
rect 50043 -5637 50053 -5585
rect 50172 -5639 50182 -5587
rect 50234 -5639 50244 -5587
rect 50364 -5638 50374 -5586
rect 50426 -5638 50436 -5586
rect 50556 -5641 50566 -5589
rect 50618 -5641 50628 -5589
rect 50750 -5640 50760 -5588
rect 50812 -5640 50822 -5588
rect 50940 -5640 50950 -5588
rect 51002 -5640 51012 -5588
rect 51135 -5638 51145 -5586
rect 51197 -5638 51207 -5586
rect 51326 -5637 51336 -5585
rect 51388 -5637 51398 -5585
rect 51521 -5639 51531 -5587
rect 51583 -5639 51593 -5587
rect 51711 -5639 51721 -5587
rect 51773 -5639 51783 -5587
rect 51901 -5638 51911 -5586
rect 51963 -5638 51973 -5586
rect 52094 -5637 52104 -5585
rect 52156 -5637 52166 -5585
rect 52285 -5637 52295 -5585
rect 52347 -5637 52357 -5585
rect 52481 -5639 52491 -5587
rect 52543 -5639 52553 -5587
rect 52670 -5639 52680 -5587
rect 52732 -5639 52742 -5587
rect 52864 -5639 52874 -5587
rect 52926 -5639 52936 -5587
rect 53053 -5639 53063 -5587
rect 53115 -5639 53125 -5587
rect 53245 -5640 53255 -5588
rect 53307 -5640 53317 -5588
rect 53438 -5640 53448 -5588
rect 53500 -5640 53510 -5588
rect 53629 -5640 53639 -5588
rect 53691 -5640 53701 -5588
rect 53821 -5639 53831 -5587
rect 53883 -5639 53893 -5587
rect 54013 -5640 54023 -5588
rect 54075 -5640 54085 -5588
rect 54206 -5640 54216 -5588
rect 54268 -5640 54278 -5588
rect 54397 -5640 54407 -5588
rect 54459 -5640 54469 -5588
rect 54589 -5639 54599 -5587
rect 54651 -5639 54661 -5587
rect 54782 -5640 54792 -5588
rect 54844 -5640 54854 -5588
rect 54974 -5640 54984 -5588
rect 55036 -5640 55046 -5588
rect 55165 -5640 55175 -5588
rect 55227 -5640 55237 -5588
rect 55356 -5640 55366 -5588
rect 55418 -5640 55428 -5588
rect 55548 -5640 55558 -5588
rect 55610 -5640 55620 -5588
rect 55741 -5639 55751 -5587
rect 55803 -5639 55813 -5587
rect 55932 -5639 55942 -5587
rect 55994 -5639 56004 -5587
rect 56126 -5640 56136 -5588
rect 56188 -5640 56198 -5588
rect 56318 -5640 56328 -5588
rect 56380 -5640 56390 -5588
rect 56510 -5640 56520 -5588
rect 56572 -5640 56582 -5588
rect 56702 -5640 56712 -5588
rect 56764 -5640 56774 -5588
rect 56894 -5640 56904 -5588
rect 56956 -5640 56966 -5588
rect 57086 -5640 57096 -5588
rect 57148 -5640 57158 -5588
rect 57278 -5640 57288 -5588
rect 57340 -5640 57350 -5588
rect 57469 -5640 57479 -5588
rect 57531 -5640 57541 -5588
rect 57661 -5640 57671 -5588
rect 57723 -5640 57733 -5588
rect 57854 -5640 57864 -5588
rect 57916 -5640 57926 -5588
rect 58046 -5640 58056 -5588
rect 58108 -5640 58118 -5588
rect 58238 -5640 58248 -5588
rect 58300 -5640 58310 -5588
rect 58429 -5640 58439 -5588
rect 58491 -5640 58501 -5588
rect 58621 -5640 58631 -5588
rect 58683 -5640 58693 -5588
rect 58812 -5640 58822 -5588
rect 58874 -5640 58884 -5588
rect 59003 -5640 59013 -5588
rect 59065 -5640 59075 -5588
rect 59197 -5640 59207 -5588
rect 59259 -5640 59269 -5588
rect 59389 -5640 59399 -5588
rect 59451 -5640 59461 -5588
rect 59582 -5639 59592 -5587
rect 59644 -5639 59654 -5587
rect 59773 -5640 59783 -5588
rect 59835 -5640 59845 -5588
rect 59965 -5640 59975 -5588
rect 60027 -5640 60037 -5588
rect 60158 -5640 60168 -5588
rect 60220 -5640 60230 -5588
rect 60350 -5640 60360 -5588
rect 60412 -5640 60422 -5588
rect 60543 -5639 60553 -5587
rect 60605 -5639 60615 -5587
rect 60734 -5640 60744 -5588
rect 60796 -5640 60806 -5588
rect 60926 -5640 60936 -5588
rect 60988 -5640 60998 -5588
rect 61117 -5640 61127 -5588
rect 61179 -5640 61189 -5588
rect 61309 -5640 61319 -5588
rect 61371 -5640 61381 -5588
rect 61501 -5640 61511 -5588
rect 61563 -5640 61573 -5588
rect 61694 -5640 61704 -5588
rect 61756 -5640 61766 -5588
rect 61885 -5640 61895 -5588
rect 61947 -5640 61957 -5588
rect 62077 -5640 62087 -5588
rect 62139 -5640 62149 -5588
rect 62269 -5639 62279 -5587
rect 62331 -5639 62341 -5587
rect 62461 -5640 62471 -5588
rect 62523 -5640 62533 -5588
rect 62651 -5640 62661 -5588
rect 62713 -5640 62723 -5588
rect 62845 -5640 62855 -5588
rect 62907 -5640 62917 -5588
rect 63037 -5639 63047 -5587
rect 63099 -5639 63109 -5587
rect 63228 -5640 63238 -5588
rect 63290 -5640 63300 -5588
rect 63421 -5640 63431 -5588
rect 63483 -5640 63493 -5588
rect 63612 -5639 63622 -5587
rect 63674 -5639 63684 -5587
rect 63804 -5640 63814 -5588
rect 63866 -5640 63876 -5588
rect 63995 -5640 64005 -5588
rect 64057 -5640 64067 -5588
rect 64189 -5639 64199 -5587
rect 64251 -5639 64261 -5587
rect 64380 -5640 64390 -5588
rect 64442 -5640 64452 -5588
rect 64572 -5640 64582 -5588
rect 64634 -5640 64644 -5588
rect 64764 -5640 64774 -5588
rect 64826 -5640 64836 -5588
rect 64956 -5640 64966 -5588
rect 65018 -5640 65028 -5588
rect 65149 -5640 65159 -5588
rect 65211 -5640 65221 -5588
rect 65340 -5640 65350 -5588
rect 65402 -5640 65412 -5588
rect 65533 -5639 65543 -5587
rect 65595 -5639 65605 -5587
rect 65724 -5640 65734 -5588
rect 65786 -5640 65796 -5588
rect 65917 -5640 65927 -5588
rect 65979 -5640 65989 -5588
rect 66108 -5640 66118 -5588
rect 66170 -5640 66180 -5588
rect 66299 -5638 66309 -5586
rect 66361 -5638 66371 -5586
rect 66494 -5640 66504 -5588
rect 66556 -5640 66566 -5588
rect 66600 -5680 66630 -5400
rect 49880 -5710 66630 -5680
rect 68000 -5710 68374 -5302
rect 51736 -5912 64284 -5878
rect 49420 -6126 49430 -6074
rect 49482 -6126 49492 -6074
rect 51736 -6382 51782 -5912
rect 52098 -6030 52146 -5912
rect 52272 -6022 52356 -5974
rect 52480 -6020 52528 -5912
rect 52654 -6024 52738 -5976
rect 52862 -6014 52910 -5912
rect 53034 -6022 53118 -5974
rect 53246 -6016 53294 -5912
rect 53424 -6022 53508 -5974
rect 53628 -6016 53676 -5912
rect 53806 -6026 53890 -5978
rect 54012 -6020 54060 -5912
rect 54190 -6026 54274 -5978
rect 54400 -6026 54448 -5912
rect 54576 -6022 54660 -5974
rect 54782 -6020 54830 -5912
rect 54960 -6026 55044 -5978
rect 55168 -6022 55216 -5912
rect 55344 -6024 55428 -5976
rect 55552 -6026 55600 -5912
rect 55726 -6022 55810 -5974
rect 55936 -6028 55984 -5912
rect 56112 -6022 56196 -5974
rect 56320 -6024 56368 -5912
rect 56494 -6022 56578 -5974
rect 56706 -6022 56754 -5912
rect 56882 -6022 56966 -5974
rect 57086 -6026 57134 -5912
rect 57260 -6018 57344 -5970
rect 57472 -6024 57520 -5912
rect 57648 -6024 57732 -5976
rect 58286 -6030 58334 -5912
rect 58464 -6022 58548 -5974
rect 58676 -6026 58724 -5912
rect 58852 -6024 58936 -5976
rect 59050 -6026 59098 -5912
rect 59234 -6030 59318 -5982
rect 59444 -6024 59492 -5912
rect 59618 -6026 59702 -5978
rect 59822 -6024 59870 -5912
rect 60002 -6026 60086 -5978
rect 60210 -6028 60258 -5912
rect 60390 -6028 60474 -5980
rect 60592 -6026 60640 -5912
rect 60774 -6022 60858 -5974
rect 60978 -6024 61026 -5912
rect 61152 -6024 61236 -5976
rect 61362 -6028 61410 -5912
rect 61538 -6026 61622 -5978
rect 61744 -6026 61792 -5912
rect 61924 -6030 62008 -5982
rect 62130 -6028 62178 -5912
rect 62308 -6028 62392 -5980
rect 62512 -6030 62560 -5912
rect 62692 -6026 62776 -5978
rect 62896 -6026 62944 -5912
rect 63076 -6024 63160 -5976
rect 63278 -6028 63326 -5912
rect 63460 -6028 63544 -5980
rect 63666 -6028 63714 -5912
rect 63846 -6028 63930 -5980
rect 51830 -6120 51910 -6114
rect 51830 -6176 51842 -6120
rect 51898 -6176 51910 -6120
rect 52037 -6123 52047 -6071
rect 52099 -6123 52109 -6071
rect 52227 -6122 52237 -6070
rect 52289 -6122 52299 -6070
rect 52419 -6121 52429 -6069
rect 52481 -6121 52491 -6069
rect 52610 -6121 52620 -6069
rect 52672 -6121 52682 -6069
rect 52804 -6121 52814 -6069
rect 52866 -6121 52876 -6069
rect 52994 -6122 53004 -6070
rect 53056 -6122 53066 -6070
rect 53188 -6121 53198 -6069
rect 53250 -6121 53260 -6069
rect 53380 -6121 53390 -6069
rect 53442 -6121 53452 -6069
rect 53571 -6122 53581 -6070
rect 53633 -6122 53643 -6070
rect 53766 -6122 53776 -6070
rect 53828 -6122 53838 -6070
rect 53956 -6122 53966 -6070
rect 54018 -6122 54028 -6070
rect 54147 -6122 54157 -6070
rect 54209 -6122 54219 -6070
rect 54339 -6122 54349 -6070
rect 54401 -6122 54411 -6070
rect 54532 -6121 54542 -6069
rect 54594 -6121 54604 -6069
rect 54724 -6122 54734 -6070
rect 54786 -6122 54796 -6070
rect 54916 -6122 54926 -6070
rect 54978 -6122 54988 -6070
rect 55109 -6122 55119 -6070
rect 55171 -6122 55181 -6070
rect 55300 -6121 55310 -6069
rect 55362 -6121 55372 -6069
rect 55492 -6122 55502 -6070
rect 55554 -6122 55564 -6070
rect 55684 -6121 55694 -6069
rect 55746 -6121 55756 -6069
rect 55876 -6121 55886 -6069
rect 55938 -6121 55948 -6069
rect 56067 -6122 56077 -6070
rect 56129 -6122 56139 -6070
rect 56260 -6121 56270 -6069
rect 56322 -6121 56332 -6069
rect 56452 -6121 56462 -6069
rect 56514 -6121 56524 -6069
rect 56646 -6122 56656 -6070
rect 56708 -6122 56718 -6070
rect 56837 -6123 56847 -6071
rect 56899 -6123 56909 -6071
rect 57026 -6122 57036 -6070
rect 57088 -6122 57098 -6070
rect 57219 -6122 57229 -6070
rect 57281 -6122 57291 -6070
rect 57412 -6122 57422 -6070
rect 57474 -6122 57484 -6070
rect 57603 -6121 57613 -6069
rect 57665 -6121 57675 -6069
rect 57794 -6121 57804 -6069
rect 57856 -6121 57866 -6069
rect 58231 -6122 58241 -6070
rect 58293 -6122 58303 -6070
rect 58421 -6121 58431 -6069
rect 58483 -6121 58493 -6069
rect 58613 -6120 58623 -6068
rect 58675 -6120 58685 -6068
rect 58804 -6120 58814 -6068
rect 58866 -6120 58876 -6068
rect 58998 -6120 59008 -6068
rect 59060 -6120 59070 -6068
rect 59188 -6121 59198 -6069
rect 59250 -6121 59260 -6069
rect 59382 -6120 59392 -6068
rect 59444 -6120 59454 -6068
rect 59574 -6120 59584 -6068
rect 59636 -6120 59646 -6068
rect 59765 -6121 59775 -6069
rect 59827 -6121 59837 -6069
rect 59960 -6121 59970 -6069
rect 60022 -6121 60032 -6069
rect 60150 -6121 60160 -6069
rect 60212 -6121 60222 -6069
rect 60341 -6121 60351 -6069
rect 60403 -6121 60413 -6069
rect 60533 -6121 60543 -6069
rect 60595 -6121 60605 -6069
rect 60726 -6120 60736 -6068
rect 60788 -6120 60798 -6068
rect 60918 -6121 60928 -6069
rect 60980 -6121 60990 -6069
rect 61110 -6121 61120 -6069
rect 61172 -6121 61182 -6069
rect 61303 -6121 61313 -6069
rect 61365 -6121 61375 -6069
rect 61494 -6120 61504 -6068
rect 61556 -6120 61566 -6068
rect 61686 -6121 61696 -6069
rect 61748 -6121 61758 -6069
rect 61878 -6120 61888 -6068
rect 61940 -6120 61950 -6068
rect 62070 -6120 62080 -6068
rect 62132 -6120 62142 -6068
rect 62261 -6121 62271 -6069
rect 62323 -6121 62333 -6069
rect 62454 -6120 62464 -6068
rect 62516 -6120 62526 -6068
rect 62646 -6120 62656 -6068
rect 62708 -6120 62718 -6068
rect 62840 -6121 62850 -6069
rect 62902 -6121 62912 -6069
rect 63031 -6122 63041 -6070
rect 63093 -6122 63103 -6070
rect 63220 -6121 63230 -6069
rect 63282 -6121 63292 -6069
rect 63413 -6121 63423 -6069
rect 63475 -6121 63485 -6069
rect 63606 -6121 63616 -6069
rect 63668 -6121 63678 -6069
rect 63797 -6120 63807 -6068
rect 63859 -6120 63869 -6068
rect 63988 -6120 63998 -6068
rect 64050 -6120 64060 -6068
rect 51830 -6182 51910 -6176
rect 64116 -6176 64196 -6170
rect 51932 -6262 51942 -6206
rect 51998 -6210 52008 -6206
rect 51998 -6262 52011 -6210
rect 52124 -6264 52134 -6208
rect 52190 -6210 52200 -6208
rect 52901 -6210 52973 -6209
rect 52190 -6262 52203 -6210
rect 52190 -6264 52200 -6262
rect 52318 -6266 52328 -6210
rect 52384 -6262 52396 -6210
rect 52384 -6266 52394 -6262
rect 52514 -6266 52524 -6210
rect 52580 -6266 52590 -6210
rect 52709 -6214 52781 -6210
rect 52704 -6270 52714 -6214
rect 52770 -6262 52781 -6214
rect 52770 -6270 52780 -6262
rect 52896 -6266 52906 -6210
rect 52962 -6261 52973 -6210
rect 53092 -6212 53164 -6210
rect 52962 -6266 52972 -6261
rect 53090 -6268 53100 -6212
rect 53156 -6268 53166 -6212
rect 53278 -6266 53288 -6210
rect 53344 -6262 53356 -6210
rect 53476 -6212 53548 -6209
rect 53344 -6266 53354 -6262
rect 53470 -6268 53480 -6212
rect 53536 -6261 53548 -6212
rect 53536 -6268 53546 -6261
rect 53662 -6264 53672 -6208
rect 53728 -6209 53738 -6208
rect 53728 -6261 53740 -6209
rect 53728 -6264 53738 -6261
rect 53860 -6266 53870 -6210
rect 53926 -6266 53936 -6210
rect 54052 -6212 54124 -6209
rect 54048 -6268 54058 -6212
rect 54114 -6268 54124 -6212
rect 54242 -6266 54252 -6210
rect 54308 -6266 54318 -6210
rect 54430 -6264 54440 -6208
rect 54496 -6209 54506 -6208
rect 54496 -6261 54507 -6209
rect 55588 -6210 55660 -6209
rect 54629 -6214 54701 -6210
rect 54819 -6212 54891 -6210
rect 55011 -6212 55083 -6210
rect 55204 -6212 55276 -6210
rect 55395 -6212 55467 -6210
rect 54496 -6264 54506 -6261
rect 54622 -6270 54632 -6214
rect 54688 -6262 54701 -6214
rect 54688 -6270 54698 -6262
rect 54816 -6268 54826 -6212
rect 54882 -6268 54892 -6212
rect 55006 -6268 55016 -6212
rect 55072 -6262 55083 -6212
rect 55072 -6268 55082 -6262
rect 55202 -6268 55212 -6212
rect 55268 -6268 55278 -6212
rect 55392 -6268 55402 -6212
rect 55458 -6268 55468 -6212
rect 55584 -6266 55594 -6210
rect 55650 -6266 55660 -6210
rect 55776 -6264 55786 -6208
rect 55842 -6210 55852 -6208
rect 55842 -6262 55853 -6210
rect 55842 -6264 55852 -6262
rect 55968 -6266 55978 -6210
rect 56034 -6266 56044 -6210
rect 56162 -6264 56172 -6208
rect 56228 -6264 56238 -6208
rect 56549 -6210 56621 -6209
rect 56355 -6212 56427 -6210
rect 56352 -6268 56362 -6212
rect 56418 -6268 56428 -6212
rect 56548 -6266 56558 -6210
rect 56614 -6266 56624 -6210
rect 56736 -6266 56746 -6210
rect 56802 -6266 56812 -6210
rect 56930 -6266 56940 -6210
rect 56996 -6266 57006 -6210
rect 57122 -6266 57132 -6210
rect 57188 -6266 57198 -6210
rect 57314 -6214 57386 -6210
rect 57507 -6212 57579 -6209
rect 57696 -6212 57768 -6209
rect 58133 -6210 58205 -6209
rect 57308 -6270 57318 -6214
rect 57374 -6262 57386 -6214
rect 57374 -6270 57384 -6262
rect 57506 -6268 57516 -6212
rect 57572 -6268 57582 -6212
rect 57692 -6268 57702 -6212
rect 57758 -6268 57768 -6212
rect 58128 -6266 58138 -6210
rect 58194 -6261 58205 -6210
rect 58325 -6212 58397 -6209
rect 58518 -6210 58590 -6209
rect 58194 -6266 58204 -6261
rect 58320 -6268 58330 -6212
rect 58386 -6261 58397 -6212
rect 58386 -6268 58396 -6261
rect 58516 -6266 58526 -6210
rect 58582 -6266 58592 -6210
rect 58710 -6212 58782 -6209
rect 58704 -6268 58714 -6212
rect 58770 -6261 58782 -6212
rect 58903 -6214 58975 -6209
rect 59095 -6212 59167 -6208
rect 58770 -6268 58780 -6261
rect 58896 -6270 58906 -6214
rect 58962 -6261 58975 -6214
rect 58962 -6270 58972 -6261
rect 59090 -6268 59100 -6212
rect 59156 -6260 59167 -6212
rect 59286 -6214 59358 -6209
rect 59478 -6212 59550 -6209
rect 59670 -6210 59742 -6208
rect 59862 -6210 59934 -6208
rect 59156 -6268 59166 -6260
rect 59282 -6270 59292 -6214
rect 59348 -6270 59358 -6214
rect 59474 -6268 59484 -6212
rect 59540 -6268 59550 -6212
rect 59668 -6266 59678 -6210
rect 59734 -6266 59744 -6210
rect 59858 -6266 59868 -6210
rect 59924 -6266 59934 -6210
rect 60054 -6214 60126 -6209
rect 60246 -6214 60318 -6208
rect 60438 -6212 60510 -6209
rect 60629 -6212 60701 -6208
rect 60050 -6270 60060 -6214
rect 60116 -6270 60126 -6214
rect 60242 -6270 60252 -6214
rect 60308 -6270 60318 -6214
rect 60434 -6268 60444 -6212
rect 60500 -6268 60510 -6212
rect 60628 -6268 60638 -6212
rect 60694 -6268 60704 -6212
rect 60823 -6214 60895 -6209
rect 61013 -6212 61085 -6209
rect 60818 -6270 60828 -6214
rect 60884 -6261 60895 -6214
rect 60884 -6270 60894 -6261
rect 61008 -6268 61018 -6212
rect 61074 -6261 61085 -6212
rect 61074 -6268 61084 -6261
rect 61202 -6264 61212 -6208
rect 61268 -6264 61278 -6208
rect 61398 -6214 61470 -6209
rect 61589 -6214 61661 -6209
rect 61782 -6214 61854 -6208
rect 61975 -6212 62047 -6209
rect 62166 -6210 62238 -6209
rect 61394 -6270 61404 -6214
rect 61460 -6270 61470 -6214
rect 61586 -6270 61596 -6214
rect 61652 -6270 61662 -6214
rect 61776 -6270 61786 -6214
rect 61842 -6260 61854 -6214
rect 61842 -6270 61852 -6260
rect 61966 -6268 61976 -6212
rect 62032 -6261 62047 -6212
rect 62032 -6268 62042 -6261
rect 62164 -6266 62174 -6210
rect 62230 -6266 62240 -6210
rect 62359 -6214 62431 -6209
rect 62549 -6212 62621 -6209
rect 62743 -6212 62815 -6208
rect 62932 -6210 63004 -6209
rect 62354 -6270 62364 -6214
rect 62420 -6261 62431 -6214
rect 62420 -6270 62430 -6261
rect 62544 -6268 62554 -6212
rect 62610 -6261 62621 -6212
rect 62610 -6268 62620 -6261
rect 62740 -6268 62750 -6212
rect 62806 -6268 62816 -6212
rect 62928 -6266 62938 -6210
rect 62994 -6266 63004 -6210
rect 63125 -6214 63197 -6209
rect 63318 -6212 63390 -6209
rect 63508 -6210 63580 -6209
rect 63124 -6270 63134 -6214
rect 63190 -6270 63200 -6214
rect 63312 -6268 63322 -6212
rect 63378 -6261 63390 -6212
rect 63378 -6268 63388 -6261
rect 63502 -6266 63512 -6210
rect 63568 -6261 63580 -6210
rect 63701 -6212 63773 -6208
rect 63890 -6210 63962 -6208
rect 63568 -6266 63578 -6261
rect 63700 -6268 63710 -6212
rect 63766 -6268 63776 -6212
rect 63890 -6260 63902 -6210
rect 63892 -6266 63902 -6260
rect 63958 -6266 63968 -6210
rect 64116 -6232 64128 -6176
rect 64184 -6232 64196 -6176
rect 64116 -6238 64196 -6232
rect 51978 -6348 52062 -6300
rect 51716 -6438 51726 -6382
rect 51782 -6422 51792 -6382
rect 52196 -6422 52244 -6302
rect 52368 -6346 52452 -6298
rect 52576 -6422 52624 -6306
rect 52754 -6348 52838 -6300
rect 52964 -6422 53012 -6310
rect 53134 -6350 53218 -6302
rect 53338 -6422 53386 -6306
rect 53520 -6350 53604 -6302
rect 53722 -6422 53770 -6300
rect 53906 -6354 53990 -6306
rect 54104 -6422 54152 -6306
rect 54290 -6352 54374 -6304
rect 54490 -6422 54538 -6306
rect 54670 -6354 54754 -6306
rect 54878 -6422 54926 -6314
rect 55056 -6352 55140 -6304
rect 55262 -6422 55310 -6306
rect 55442 -6356 55526 -6308
rect 55652 -6422 55700 -6302
rect 55824 -6360 55908 -6312
rect 56028 -6422 56076 -6314
rect 56210 -6366 56294 -6318
rect 56410 -6422 56458 -6314
rect 56590 -6352 56674 -6304
rect 56796 -6422 56844 -6314
rect 56976 -6346 57060 -6298
rect 57188 -6422 57236 -6310
rect 57360 -6358 57444 -6310
rect 57568 -6422 57616 -6304
rect 57746 -6352 57830 -6304
rect 58178 -6358 58262 -6310
rect 58382 -6422 58430 -6306
rect 58564 -6358 58648 -6310
rect 58774 -6422 58822 -6310
rect 58946 -6352 59030 -6304
rect 59150 -6422 59198 -6304
rect 59330 -6358 59414 -6310
rect 59542 -6422 59590 -6308
rect 59716 -6358 59800 -6310
rect 59914 -6422 59962 -6310
rect 60098 -6352 60182 -6304
rect 60306 -6422 60354 -6310
rect 60486 -6350 60570 -6302
rect 60688 -6422 60736 -6304
rect 60868 -6346 60952 -6298
rect 61074 -6422 61122 -6310
rect 61252 -6350 61336 -6302
rect 61460 -6422 61508 -6304
rect 61634 -6352 61718 -6304
rect 61842 -6422 61890 -6304
rect 62018 -6350 62102 -6302
rect 62218 -6422 62266 -6304
rect 62404 -6346 62488 -6298
rect 62610 -6422 62658 -6306
rect 62786 -6348 62870 -6300
rect 62994 -6422 63042 -6308
rect 63172 -6346 63256 -6298
rect 63384 -6422 63432 -6306
rect 63554 -6346 63638 -6298
rect 63760 -6422 63808 -6302
rect 63940 -6348 64024 -6300
rect 64230 -6400 64284 -5912
rect 66908 -6002 66918 -5950
rect 66970 -6002 66980 -5950
rect 68000 -6298 68362 -5710
rect 68920 -6272 68930 -5188
rect 69296 -6272 69306 -5188
rect 64226 -6422 64236 -6400
rect 51782 -6438 64236 -6422
rect 51736 -6456 64236 -6438
rect 64292 -6456 64302 -6400
rect 51846 -6570 64140 -6542
rect 47244 -7752 47254 -6678
rect 47614 -7752 47624 -6678
rect 48194 -7240 48556 -6644
rect 49426 -6924 49436 -6872
rect 49488 -6924 49498 -6872
rect 51846 -6996 51884 -6570
rect 52096 -6650 52154 -6570
rect 52272 -6646 52378 -6616
rect 52482 -6646 52540 -6570
rect 52652 -6646 52758 -6616
rect 52864 -6638 52920 -6570
rect 53034 -6640 53140 -6610
rect 53250 -6630 53298 -6570
rect 53406 -6636 53512 -6606
rect 53642 -6628 53686 -6570
rect 53800 -6642 53906 -6612
rect 54020 -6634 54066 -6570
rect 54182 -6640 54288 -6610
rect 54404 -6624 54460 -6570
rect 54570 -6642 54676 -6612
rect 54790 -6628 54838 -6570
rect 54954 -6646 55060 -6616
rect 55168 -6630 55220 -6570
rect 55340 -6648 55446 -6618
rect 55554 -6630 55610 -6570
rect 55714 -6646 55820 -6616
rect 55940 -6636 55992 -6570
rect 56096 -6646 56202 -6616
rect 56322 -6634 56376 -6570
rect 56474 -6644 56580 -6614
rect 56708 -6632 56760 -6570
rect 56874 -6638 56980 -6608
rect 57088 -6632 57148 -6570
rect 57248 -6640 57354 -6610
rect 57476 -6636 57522 -6570
rect 57646 -6648 57752 -6618
rect 58280 -6622 58338 -6570
rect 58452 -6640 58558 -6610
rect 58664 -6622 58720 -6570
rect 58836 -6638 58942 -6608
rect 59044 -6614 59108 -6570
rect 59216 -6638 59322 -6608
rect 59444 -6620 59478 -6570
rect 59596 -6632 59702 -6602
rect 59818 -6622 59872 -6570
rect 59974 -6636 60080 -6606
rect 60202 -6620 60252 -6570
rect 60360 -6646 60466 -6616
rect 60584 -6618 60640 -6570
rect 60754 -6634 60860 -6604
rect 60972 -6630 61024 -6570
rect 61132 -6634 61238 -6604
rect 61352 -6632 61404 -6570
rect 61526 -6636 61632 -6606
rect 61736 -6628 61788 -6570
rect 61916 -6638 62022 -6608
rect 62124 -6640 62176 -6570
rect 62286 -6634 62392 -6604
rect 62504 -6632 62556 -6570
rect 62676 -6638 62782 -6608
rect 62888 -6634 62940 -6570
rect 63058 -6634 63164 -6604
rect 63274 -6636 63326 -6570
rect 63446 -6638 63552 -6608
rect 63656 -6638 63708 -6570
rect 63830 -6638 63936 -6608
rect 52038 -6690 52110 -6689
rect 52034 -6746 52044 -6690
rect 52100 -6746 52110 -6690
rect 52228 -6690 52300 -6688
rect 52228 -6746 52238 -6690
rect 52294 -6746 52304 -6690
rect 52420 -6696 52492 -6687
rect 52611 -6692 52683 -6687
rect 52805 -6692 52877 -6687
rect 52995 -6692 53067 -6688
rect 53189 -6690 53261 -6687
rect 53381 -6690 53453 -6687
rect 52420 -6739 52432 -6696
rect 52422 -6752 52432 -6739
rect 52488 -6752 52498 -6696
rect 52611 -6739 52622 -6692
rect 52612 -6748 52622 -6739
rect 52678 -6748 52688 -6692
rect 52805 -6739 52818 -6692
rect 52808 -6748 52818 -6739
rect 52874 -6748 52884 -6692
rect 52995 -6740 53006 -6692
rect 52996 -6748 53006 -6740
rect 53062 -6748 53072 -6692
rect 53189 -6739 53200 -6690
rect 53190 -6746 53200 -6739
rect 53256 -6746 53266 -6690
rect 53381 -6739 53394 -6690
rect 53384 -6746 53394 -6739
rect 53450 -6746 53460 -6690
rect 53572 -6692 53644 -6688
rect 53767 -6690 53839 -6688
rect 53572 -6748 53582 -6692
rect 53638 -6748 53648 -6692
rect 53764 -6746 53774 -6690
rect 53830 -6746 53840 -6690
rect 53957 -6694 54029 -6688
rect 54148 -6692 54220 -6688
rect 53954 -6750 53964 -6694
rect 54020 -6750 54030 -6694
rect 54146 -6748 54156 -6692
rect 54212 -6748 54222 -6692
rect 54340 -6694 54412 -6688
rect 54533 -6690 54605 -6687
rect 54340 -6750 54350 -6694
rect 54406 -6750 54416 -6694
rect 54532 -6746 54542 -6690
rect 54598 -6746 54608 -6690
rect 54725 -6692 54797 -6688
rect 54917 -6690 54989 -6688
rect 54725 -6740 54740 -6692
rect 54730 -6748 54740 -6740
rect 54796 -6748 54806 -6692
rect 54916 -6746 54926 -6690
rect 54982 -6746 54992 -6690
rect 55110 -6696 55182 -6688
rect 55301 -6692 55373 -6687
rect 55110 -6752 55120 -6696
rect 55176 -6752 55186 -6696
rect 55300 -6748 55310 -6692
rect 55366 -6748 55376 -6692
rect 55493 -6696 55565 -6688
rect 55685 -6690 55757 -6687
rect 55492 -6752 55502 -6696
rect 55558 -6752 55568 -6696
rect 55680 -6746 55690 -6690
rect 55746 -6739 55757 -6690
rect 55877 -6694 55949 -6687
rect 55746 -6746 55756 -6739
rect 55876 -6750 55886 -6694
rect 55942 -6750 55952 -6694
rect 56068 -6744 56078 -6688
rect 56134 -6744 56144 -6688
rect 56261 -6692 56333 -6687
rect 56261 -6739 56272 -6692
rect 56262 -6748 56272 -6739
rect 56328 -6748 56338 -6692
rect 56453 -6694 56525 -6687
rect 56647 -6694 56719 -6688
rect 56838 -6690 56910 -6689
rect 56450 -6750 56460 -6694
rect 56516 -6750 56526 -6694
rect 56647 -6740 56658 -6694
rect 56648 -6750 56658 -6740
rect 56714 -6750 56724 -6694
rect 56838 -6746 56848 -6690
rect 56904 -6746 56914 -6690
rect 57027 -6696 57099 -6688
rect 57220 -6690 57292 -6688
rect 57027 -6740 57038 -6696
rect 57028 -6752 57038 -6740
rect 57094 -6752 57104 -6696
rect 57218 -6746 57228 -6690
rect 57284 -6746 57294 -6690
rect 57413 -6696 57485 -6688
rect 57604 -6692 57676 -6687
rect 57412 -6752 57422 -6696
rect 57478 -6752 57488 -6696
rect 57598 -6748 57608 -6692
rect 57664 -6739 57676 -6692
rect 57795 -6694 57867 -6687
rect 58226 -6694 58298 -6688
rect 58416 -6692 58488 -6687
rect 57795 -6739 57806 -6694
rect 57664 -6748 57674 -6739
rect 57796 -6750 57806 -6739
rect 57862 -6750 57872 -6694
rect 58220 -6750 58230 -6694
rect 58286 -6740 58298 -6694
rect 58286 -6750 58296 -6740
rect 58410 -6748 58420 -6692
rect 58476 -6739 58488 -6692
rect 58608 -6698 58680 -6686
rect 58799 -6692 58871 -6686
rect 58476 -6748 58486 -6739
rect 58602 -6754 58612 -6698
rect 58668 -6738 58680 -6698
rect 58668 -6754 58678 -6738
rect 58792 -6748 58802 -6692
rect 58858 -6738 58871 -6692
rect 58993 -6694 59065 -6686
rect 59183 -6690 59255 -6687
rect 58858 -6748 58868 -6738
rect 58986 -6750 58996 -6694
rect 59052 -6738 59065 -6694
rect 59052 -6750 59062 -6738
rect 59180 -6746 59190 -6690
rect 59246 -6746 59256 -6690
rect 59377 -6694 59449 -6686
rect 59569 -6692 59641 -6686
rect 59372 -6750 59382 -6694
rect 59438 -6738 59449 -6694
rect 59438 -6750 59448 -6738
rect 59562 -6748 59572 -6692
rect 59628 -6738 59641 -6692
rect 59760 -6694 59832 -6687
rect 59955 -6690 60027 -6687
rect 59628 -6748 59638 -6738
rect 59754 -6750 59764 -6694
rect 59820 -6739 59832 -6694
rect 59820 -6750 59830 -6739
rect 59950 -6746 59960 -6690
rect 60016 -6739 60027 -6690
rect 60145 -6692 60217 -6687
rect 60336 -6690 60408 -6687
rect 60016 -6746 60026 -6739
rect 60144 -6748 60154 -6692
rect 60210 -6748 60220 -6692
rect 60332 -6746 60342 -6690
rect 60398 -6746 60408 -6690
rect 60528 -6696 60600 -6687
rect 60721 -6688 60793 -6686
rect 60524 -6752 60534 -6696
rect 60590 -6752 60600 -6696
rect 60716 -6744 60726 -6688
rect 60782 -6738 60793 -6688
rect 60913 -6694 60985 -6687
rect 61105 -6690 61177 -6687
rect 60782 -6744 60792 -6738
rect 60908 -6750 60918 -6694
rect 60974 -6739 60985 -6694
rect 60974 -6750 60984 -6739
rect 61100 -6746 61110 -6690
rect 61166 -6739 61177 -6690
rect 61298 -6694 61370 -6687
rect 61489 -6690 61561 -6686
rect 61166 -6746 61176 -6739
rect 61290 -6750 61300 -6694
rect 61356 -6739 61370 -6694
rect 61356 -6750 61366 -6739
rect 61482 -6746 61492 -6690
rect 61548 -6738 61561 -6690
rect 61681 -6696 61753 -6687
rect 61873 -6690 61945 -6686
rect 61548 -6746 61558 -6738
rect 61678 -6752 61688 -6696
rect 61744 -6752 61754 -6696
rect 61864 -6746 61874 -6690
rect 61930 -6738 61945 -6690
rect 62065 -6692 62137 -6686
rect 62256 -6690 62328 -6687
rect 61930 -6746 61940 -6738
rect 62060 -6748 62070 -6692
rect 62126 -6738 62137 -6692
rect 62126 -6748 62136 -6738
rect 62250 -6746 62260 -6690
rect 62316 -6739 62328 -6690
rect 62449 -6692 62521 -6686
rect 62641 -6690 62713 -6686
rect 62835 -6690 62907 -6687
rect 62316 -6746 62326 -6739
rect 62446 -6748 62456 -6692
rect 62512 -6748 62522 -6692
rect 62634 -6746 62644 -6690
rect 62700 -6738 62713 -6690
rect 62700 -6746 62710 -6738
rect 62830 -6746 62840 -6690
rect 62896 -6739 62907 -6690
rect 63026 -6692 63098 -6688
rect 63215 -6692 63287 -6687
rect 63408 -6692 63480 -6687
rect 63601 -6690 63673 -6687
rect 63792 -6688 63864 -6686
rect 62896 -6746 62906 -6739
rect 63018 -6748 63028 -6692
rect 63084 -6740 63098 -6692
rect 63084 -6748 63094 -6740
rect 63210 -6748 63220 -6692
rect 63276 -6739 63287 -6692
rect 63276 -6748 63286 -6739
rect 63402 -6748 63412 -6692
rect 63468 -6739 63480 -6692
rect 63468 -6748 63478 -6739
rect 63598 -6746 63608 -6690
rect 63664 -6746 63674 -6690
rect 63786 -6744 63796 -6688
rect 63852 -6738 63864 -6688
rect 63983 -6690 64055 -6686
rect 63852 -6744 63862 -6738
rect 63982 -6746 63992 -6690
rect 64048 -6746 64058 -6690
rect 51940 -6880 51950 -6828
rect 52002 -6880 52012 -6828
rect 52132 -6880 52142 -6828
rect 52194 -6880 52204 -6828
rect 52325 -6880 52335 -6828
rect 52387 -6880 52397 -6828
rect 52517 -6880 52527 -6828
rect 52579 -6880 52589 -6828
rect 52710 -6880 52720 -6828
rect 52772 -6880 52782 -6828
rect 52902 -6879 52912 -6827
rect 52964 -6879 52974 -6827
rect 53093 -6880 53103 -6828
rect 53155 -6880 53165 -6828
rect 53285 -6880 53295 -6828
rect 53347 -6880 53357 -6828
rect 53477 -6879 53487 -6827
rect 53539 -6879 53549 -6827
rect 53669 -6879 53679 -6827
rect 53731 -6879 53741 -6827
rect 53861 -6880 53871 -6828
rect 53923 -6880 53933 -6828
rect 54053 -6879 54063 -6827
rect 54115 -6879 54125 -6827
rect 54245 -6880 54255 -6828
rect 54307 -6880 54317 -6828
rect 54436 -6879 54446 -6827
rect 54498 -6879 54508 -6827
rect 54630 -6880 54640 -6828
rect 54692 -6880 54702 -6828
rect 54820 -6880 54830 -6828
rect 54882 -6880 54892 -6828
rect 55012 -6880 55022 -6828
rect 55074 -6880 55084 -6828
rect 55205 -6880 55215 -6828
rect 55267 -6880 55277 -6828
rect 55396 -6880 55406 -6828
rect 55458 -6880 55468 -6828
rect 55589 -6879 55599 -6827
rect 55651 -6879 55661 -6827
rect 55782 -6880 55792 -6828
rect 55844 -6880 55854 -6828
rect 55973 -6880 55983 -6828
rect 56035 -6880 56045 -6828
rect 56166 -6880 56176 -6828
rect 56228 -6880 56238 -6828
rect 56356 -6880 56366 -6828
rect 56418 -6880 56428 -6828
rect 56550 -6879 56560 -6827
rect 56612 -6879 56622 -6827
rect 56739 -6880 56749 -6828
rect 56801 -6880 56811 -6828
rect 56932 -6880 56942 -6828
rect 56994 -6880 57004 -6828
rect 57125 -6880 57135 -6828
rect 57187 -6880 57197 -6828
rect 57315 -6880 57325 -6828
rect 57377 -6880 57387 -6828
rect 57508 -6879 57518 -6827
rect 57570 -6879 57580 -6827
rect 57697 -6879 57707 -6827
rect 57759 -6879 57769 -6827
rect 58130 -6879 58138 -6827
rect 58190 -6879 58200 -6827
rect 58320 -6879 58330 -6827
rect 58382 -6879 58392 -6827
rect 58513 -6879 58523 -6827
rect 58575 -6879 58585 -6827
rect 58705 -6879 58715 -6827
rect 58767 -6879 58777 -6827
rect 58898 -6879 58908 -6827
rect 58960 -6879 58970 -6827
rect 59090 -6878 59100 -6826
rect 59152 -6878 59162 -6826
rect 59281 -6879 59291 -6827
rect 59343 -6879 59353 -6827
rect 59473 -6879 59483 -6827
rect 59535 -6879 59545 -6827
rect 59665 -6878 59675 -6826
rect 59727 -6878 59737 -6826
rect 59857 -6878 59867 -6826
rect 59919 -6878 59929 -6826
rect 60049 -6879 60059 -6827
rect 60111 -6879 60121 -6827
rect 60241 -6878 60251 -6826
rect 60303 -6878 60313 -6826
rect 60433 -6879 60443 -6827
rect 60495 -6879 60505 -6827
rect 60624 -6878 60634 -6826
rect 60686 -6878 60696 -6826
rect 60818 -6879 60828 -6827
rect 60880 -6879 60890 -6827
rect 61008 -6879 61018 -6827
rect 61070 -6879 61080 -6827
rect 61200 -6879 61210 -6827
rect 61262 -6879 61272 -6827
rect 61393 -6879 61403 -6827
rect 61455 -6879 61465 -6827
rect 61584 -6879 61594 -6827
rect 61646 -6879 61656 -6827
rect 61777 -6878 61787 -6826
rect 61839 -6878 61849 -6826
rect 61970 -6879 61980 -6827
rect 62032 -6879 62042 -6827
rect 62161 -6879 62171 -6827
rect 62223 -6879 62233 -6827
rect 62354 -6879 62364 -6827
rect 62416 -6879 62426 -6827
rect 62544 -6879 62554 -6827
rect 62606 -6879 62616 -6827
rect 62738 -6878 62748 -6826
rect 62800 -6878 62810 -6826
rect 62927 -6879 62937 -6827
rect 62989 -6879 62999 -6827
rect 63120 -6879 63130 -6827
rect 63182 -6879 63192 -6827
rect 63313 -6879 63323 -6827
rect 63375 -6879 63385 -6827
rect 63503 -6879 63513 -6827
rect 63565 -6879 63575 -6827
rect 63696 -6878 63706 -6826
rect 63758 -6878 63768 -6826
rect 63885 -6878 63895 -6826
rect 63947 -6878 63957 -6826
rect 51998 -6996 52058 -6926
rect 52162 -6958 52268 -6928
rect 52382 -6996 52438 -6928
rect 52554 -6960 52660 -6930
rect 52762 -6996 52826 -6928
rect 52936 -6954 53042 -6924
rect 53150 -6996 53204 -6934
rect 53312 -6966 53418 -6936
rect 53538 -6996 53584 -6934
rect 53698 -6964 53804 -6934
rect 53922 -6996 53966 -6938
rect 54092 -6962 54198 -6932
rect 54304 -6996 54352 -6942
rect 54482 -6954 54588 -6924
rect 54688 -6996 54738 -6942
rect 54848 -6960 54954 -6930
rect 55072 -6996 55122 -6938
rect 55238 -6960 55344 -6930
rect 55452 -6996 55508 -6938
rect 55636 -6958 55742 -6928
rect 55838 -6996 55890 -6940
rect 56008 -6968 56114 -6938
rect 56226 -6996 56270 -6936
rect 56394 -6966 56500 -6936
rect 56608 -6996 56660 -6938
rect 56772 -6960 56878 -6930
rect 56992 -6996 57040 -6938
rect 57168 -6962 57274 -6932
rect 57374 -6996 57424 -6936
rect 57546 -6968 57652 -6938
rect 57756 -6996 57810 -6942
rect 58174 -6996 58230 -6928
rect 58340 -6952 58446 -6922
rect 58560 -6996 58614 -6928
rect 58744 -6954 58850 -6924
rect 58948 -6996 58994 -6930
rect 59130 -6950 59236 -6920
rect 59340 -6996 59378 -6932
rect 59512 -6950 59618 -6920
rect 59716 -6996 59768 -6930
rect 59892 -6950 59998 -6920
rect 60104 -6996 60146 -6932
rect 60282 -6960 60388 -6930
rect 60480 -6996 60532 -6932
rect 60662 -6960 60768 -6930
rect 60868 -6996 60920 -6928
rect 61042 -6952 61148 -6922
rect 61254 -6996 61306 -6932
rect 61420 -6956 61526 -6926
rect 61638 -6996 61690 -6928
rect 61808 -6952 61914 -6922
rect 62028 -6996 62080 -6930
rect 62206 -6960 62312 -6930
rect 62410 -6996 62462 -6934
rect 62580 -6960 62686 -6930
rect 62798 -6996 62850 -6932
rect 62964 -6950 63070 -6920
rect 63174 -6996 63226 -6934
rect 63348 -6956 63454 -6926
rect 63562 -6996 63614 -6932
rect 63732 -6954 63838 -6924
rect 63940 -6996 63992 -6934
rect 64112 -6996 64140 -6570
rect 66902 -6902 66912 -6850
rect 66964 -6902 66974 -6850
rect 51846 -7024 64140 -6996
rect 48190 -7640 48556 -7240
rect 49890 -7260 66624 -7230
rect 49890 -7540 49920 -7260
rect 50077 -7354 50087 -7302
rect 50139 -7354 50149 -7302
rect 50267 -7353 50277 -7301
rect 50329 -7353 50339 -7301
rect 50460 -7356 50470 -7304
rect 50522 -7356 50532 -7304
rect 50652 -7351 50662 -7299
rect 50714 -7351 50724 -7299
rect 50844 -7355 50854 -7303
rect 50906 -7355 50916 -7303
rect 51036 -7350 51046 -7298
rect 51098 -7350 51108 -7298
rect 51228 -7351 51238 -7299
rect 51290 -7351 51300 -7299
rect 51418 -7350 51428 -7298
rect 51480 -7350 51490 -7298
rect 51612 -7361 51622 -7309
rect 51674 -7361 51684 -7309
rect 51801 -7359 51811 -7307
rect 51863 -7359 51873 -7307
rect 51991 -7359 52001 -7307
rect 52053 -7359 52063 -7307
rect 52190 -7360 52200 -7308
rect 52252 -7360 52262 -7308
rect 52382 -7359 52392 -7307
rect 52444 -7359 52454 -7307
rect 52572 -7360 52582 -7308
rect 52634 -7360 52644 -7308
rect 52764 -7353 52774 -7301
rect 52826 -7353 52836 -7301
rect 52956 -7303 53028 -7298
rect 52956 -7355 52966 -7303
rect 53018 -7355 53028 -7303
rect 53149 -7354 53159 -7302
rect 53211 -7354 53221 -7302
rect 53341 -7352 53351 -7300
rect 53403 -7352 53413 -7300
rect 53532 -7352 53542 -7300
rect 53594 -7352 53604 -7300
rect 53726 -7357 53736 -7305
rect 53788 -7357 53798 -7305
rect 53917 -7353 53927 -7301
rect 53979 -7353 53989 -7301
rect 54109 -7349 54119 -7297
rect 54171 -7349 54181 -7297
rect 54302 -7353 54312 -7301
rect 54364 -7353 54374 -7301
rect 54494 -7353 54504 -7301
rect 54556 -7353 54566 -7301
rect 54687 -7354 54697 -7302
rect 54749 -7354 54759 -7302
rect 54879 -7352 54889 -7300
rect 54941 -7352 54951 -7300
rect 55070 -7351 55080 -7299
rect 55132 -7351 55142 -7299
rect 55261 -7350 55271 -7298
rect 55323 -7350 55333 -7298
rect 55454 -7350 55464 -7298
rect 55516 -7350 55526 -7298
rect 55645 -7359 55655 -7307
rect 55707 -7359 55717 -7307
rect 55836 -7360 55846 -7308
rect 55898 -7360 55908 -7308
rect 56026 -7361 56036 -7309
rect 56088 -7361 56098 -7309
rect 56220 -7365 56230 -7313
rect 56282 -7365 56292 -7313
rect 56412 -7367 56422 -7315
rect 56474 -7367 56484 -7315
rect 56606 -7366 56616 -7314
rect 56668 -7366 56678 -7314
rect 56798 -7363 56808 -7311
rect 56860 -7363 56870 -7311
rect 56987 -7360 56997 -7308
rect 57049 -7360 57059 -7308
rect 57181 -7358 57191 -7306
rect 57243 -7358 57253 -7306
rect 57374 -7359 57384 -7307
rect 57436 -7359 57446 -7307
rect 57567 -7360 57577 -7308
rect 57629 -7360 57639 -7308
rect 57756 -7360 57766 -7308
rect 57818 -7360 57828 -7308
rect 57949 -7360 57959 -7308
rect 58011 -7360 58021 -7308
rect 58141 -7360 58151 -7308
rect 58203 -7360 58213 -7308
rect 58332 -7360 58342 -7308
rect 58394 -7360 58404 -7308
rect 58525 -7360 58535 -7308
rect 58587 -7360 58597 -7308
rect 58716 -7359 58726 -7307
rect 58778 -7359 58788 -7307
rect 58911 -7360 58921 -7308
rect 58973 -7360 58983 -7308
rect 59100 -7360 59110 -7308
rect 59162 -7360 59172 -7308
rect 59293 -7360 59303 -7308
rect 59355 -7360 59365 -7308
rect 59485 -7360 59495 -7308
rect 59547 -7360 59557 -7308
rect 59676 -7360 59686 -7308
rect 59738 -7360 59748 -7308
rect 59868 -7360 59878 -7308
rect 59930 -7360 59940 -7308
rect 60061 -7360 60071 -7308
rect 60123 -7360 60133 -7308
rect 60250 -7361 60260 -7309
rect 60312 -7361 60322 -7309
rect 60444 -7360 60454 -7308
rect 60506 -7360 60516 -7308
rect 60635 -7360 60645 -7308
rect 60697 -7360 60707 -7308
rect 60828 -7360 60838 -7308
rect 60890 -7360 60900 -7308
rect 61020 -7360 61030 -7308
rect 61082 -7360 61092 -7308
rect 61212 -7361 61222 -7309
rect 61274 -7361 61284 -7309
rect 61405 -7359 61415 -7307
rect 61467 -7359 61477 -7307
rect 61595 -7359 61605 -7307
rect 61657 -7359 61667 -7307
rect 61788 -7361 61798 -7309
rect 61850 -7361 61860 -7309
rect 61980 -7360 61990 -7308
rect 62042 -7360 62052 -7308
rect 62173 -7359 62183 -7307
rect 62235 -7359 62245 -7307
rect 62364 -7359 62374 -7307
rect 62426 -7359 62436 -7307
rect 62556 -7360 62566 -7308
rect 62618 -7360 62628 -7308
rect 62747 -7360 62757 -7308
rect 62809 -7360 62819 -7308
rect 62939 -7360 62949 -7308
rect 63001 -7360 63011 -7308
rect 63133 -7359 63143 -7307
rect 63195 -7359 63205 -7307
rect 63325 -7360 63335 -7308
rect 63387 -7360 63397 -7308
rect 63515 -7361 63525 -7309
rect 63577 -7361 63587 -7309
rect 63706 -7362 63716 -7310
rect 63768 -7362 63778 -7310
rect 63899 -7360 63909 -7308
rect 63961 -7360 63971 -7308
rect 64092 -7359 64102 -7307
rect 64154 -7359 64164 -7307
rect 64285 -7360 64295 -7308
rect 64347 -7360 64357 -7308
rect 64476 -7360 64486 -7308
rect 64538 -7360 64548 -7308
rect 64667 -7360 64677 -7308
rect 64729 -7360 64739 -7308
rect 64860 -7360 64870 -7308
rect 64922 -7360 64932 -7308
rect 65053 -7360 65063 -7308
rect 65115 -7360 65125 -7308
rect 65244 -7360 65254 -7308
rect 65306 -7360 65316 -7308
rect 65435 -7359 65445 -7307
rect 65497 -7359 65507 -7307
rect 65626 -7359 65636 -7307
rect 65688 -7359 65698 -7307
rect 65819 -7360 65829 -7308
rect 65881 -7360 65891 -7308
rect 66013 -7360 66023 -7308
rect 66075 -7360 66085 -7308
rect 66201 -7361 66211 -7309
rect 66263 -7361 66273 -7309
rect 66395 -7369 66405 -7317
rect 66457 -7369 66467 -7317
rect 49981 -7497 49991 -7445
rect 50043 -7497 50053 -7445
rect 50172 -7499 50182 -7447
rect 50234 -7499 50244 -7447
rect 50364 -7498 50374 -7446
rect 50426 -7498 50436 -7446
rect 50556 -7501 50566 -7449
rect 50618 -7501 50628 -7449
rect 50750 -7500 50760 -7448
rect 50812 -7500 50822 -7448
rect 50940 -7500 50950 -7448
rect 51002 -7500 51012 -7448
rect 51135 -7498 51145 -7446
rect 51197 -7498 51207 -7446
rect 51326 -7497 51336 -7445
rect 51388 -7497 51398 -7445
rect 51521 -7499 51531 -7447
rect 51583 -7499 51593 -7447
rect 51711 -7499 51721 -7447
rect 51773 -7499 51783 -7447
rect 51901 -7498 51911 -7446
rect 51963 -7498 51973 -7446
rect 52094 -7497 52104 -7445
rect 52156 -7497 52166 -7445
rect 52285 -7497 52295 -7445
rect 52347 -7497 52357 -7445
rect 52481 -7499 52491 -7447
rect 52543 -7499 52553 -7447
rect 52670 -7499 52680 -7447
rect 52732 -7499 52742 -7447
rect 52864 -7499 52874 -7447
rect 52926 -7499 52936 -7447
rect 53053 -7499 53063 -7447
rect 53115 -7499 53125 -7447
rect 53245 -7500 53255 -7448
rect 53307 -7500 53317 -7448
rect 53438 -7500 53448 -7448
rect 53500 -7500 53510 -7448
rect 53629 -7500 53639 -7448
rect 53691 -7500 53701 -7448
rect 53821 -7499 53831 -7447
rect 53883 -7499 53893 -7447
rect 54013 -7500 54023 -7448
rect 54075 -7500 54085 -7448
rect 54206 -7500 54216 -7448
rect 54268 -7500 54278 -7448
rect 54397 -7500 54407 -7448
rect 54459 -7500 54469 -7448
rect 54589 -7499 54599 -7447
rect 54651 -7499 54661 -7447
rect 54782 -7500 54792 -7448
rect 54844 -7500 54854 -7448
rect 54974 -7500 54984 -7448
rect 55036 -7500 55046 -7448
rect 55165 -7500 55175 -7448
rect 55227 -7500 55237 -7448
rect 55356 -7500 55366 -7448
rect 55418 -7500 55428 -7448
rect 55548 -7500 55558 -7448
rect 55610 -7500 55620 -7448
rect 55741 -7499 55751 -7447
rect 55803 -7499 55813 -7447
rect 55932 -7499 55942 -7447
rect 55994 -7499 56004 -7447
rect 56126 -7500 56136 -7448
rect 56188 -7500 56198 -7448
rect 56318 -7500 56328 -7448
rect 56380 -7500 56390 -7448
rect 56510 -7500 56520 -7448
rect 56572 -7500 56582 -7448
rect 56702 -7500 56712 -7448
rect 56764 -7500 56774 -7448
rect 56894 -7500 56904 -7448
rect 56956 -7500 56966 -7448
rect 57086 -7500 57096 -7448
rect 57148 -7500 57158 -7448
rect 57278 -7500 57288 -7448
rect 57340 -7500 57350 -7448
rect 57469 -7500 57479 -7448
rect 57531 -7500 57541 -7448
rect 57661 -7500 57671 -7448
rect 57723 -7500 57733 -7448
rect 57854 -7500 57864 -7448
rect 57916 -7500 57926 -7448
rect 58046 -7500 58056 -7448
rect 58108 -7500 58118 -7448
rect 58238 -7500 58248 -7448
rect 58300 -7500 58310 -7448
rect 58429 -7500 58439 -7448
rect 58491 -7500 58501 -7448
rect 58621 -7500 58631 -7448
rect 58683 -7500 58693 -7448
rect 58812 -7500 58822 -7448
rect 58874 -7500 58884 -7448
rect 59003 -7500 59013 -7448
rect 59065 -7500 59075 -7448
rect 59197 -7500 59207 -7448
rect 59259 -7500 59269 -7448
rect 59389 -7500 59399 -7448
rect 59451 -7500 59461 -7448
rect 59582 -7499 59592 -7447
rect 59644 -7499 59654 -7447
rect 59773 -7500 59783 -7448
rect 59835 -7500 59845 -7448
rect 59965 -7500 59975 -7448
rect 60027 -7500 60037 -7448
rect 60158 -7500 60168 -7448
rect 60220 -7500 60230 -7448
rect 60350 -7500 60360 -7448
rect 60412 -7500 60422 -7448
rect 60543 -7499 60553 -7447
rect 60605 -7499 60615 -7447
rect 60734 -7500 60744 -7448
rect 60796 -7500 60806 -7448
rect 60926 -7500 60936 -7448
rect 60988 -7500 60998 -7448
rect 61117 -7500 61127 -7448
rect 61179 -7500 61189 -7448
rect 61309 -7500 61319 -7448
rect 61371 -7500 61381 -7448
rect 61501 -7500 61511 -7448
rect 61563 -7500 61573 -7448
rect 61694 -7500 61704 -7448
rect 61756 -7500 61766 -7448
rect 61885 -7500 61895 -7448
rect 61947 -7500 61957 -7448
rect 62077 -7500 62087 -7448
rect 62139 -7500 62149 -7448
rect 62269 -7499 62279 -7447
rect 62331 -7499 62341 -7447
rect 62461 -7500 62471 -7448
rect 62523 -7500 62533 -7448
rect 62651 -7500 62661 -7448
rect 62713 -7500 62723 -7448
rect 62845 -7500 62855 -7448
rect 62907 -7500 62917 -7448
rect 63037 -7499 63047 -7447
rect 63099 -7499 63109 -7447
rect 63228 -7500 63238 -7448
rect 63290 -7500 63300 -7448
rect 63421 -7500 63431 -7448
rect 63483 -7500 63493 -7448
rect 63612 -7499 63622 -7447
rect 63674 -7499 63684 -7447
rect 63804 -7500 63814 -7448
rect 63866 -7500 63876 -7448
rect 63995 -7500 64005 -7448
rect 64057 -7500 64067 -7448
rect 64189 -7499 64199 -7447
rect 64251 -7499 64261 -7447
rect 64380 -7500 64390 -7448
rect 64442 -7500 64452 -7448
rect 64572 -7500 64582 -7448
rect 64634 -7500 64644 -7448
rect 64764 -7500 64774 -7448
rect 64826 -7500 64836 -7448
rect 64956 -7500 64966 -7448
rect 65018 -7500 65028 -7448
rect 65149 -7500 65159 -7448
rect 65211 -7500 65221 -7448
rect 65340 -7500 65350 -7448
rect 65402 -7500 65412 -7448
rect 65533 -7499 65543 -7447
rect 65595 -7499 65605 -7447
rect 65724 -7500 65734 -7448
rect 65786 -7500 65796 -7448
rect 65917 -7500 65927 -7448
rect 65979 -7500 65989 -7448
rect 66108 -7500 66118 -7448
rect 66170 -7500 66180 -7448
rect 66299 -7498 66309 -7446
rect 66361 -7498 66371 -7446
rect 66494 -7500 66504 -7448
rect 66556 -7500 66566 -7448
rect 66594 -7540 66624 -7260
rect 49890 -7570 66624 -7540
rect 68006 -7234 68368 -6644
rect 68006 -7640 68374 -7234
rect 68368 -7642 68374 -7640
rect 49928 -7664 66600 -7658
rect 48262 -7706 48458 -7700
rect 48262 -7764 48274 -7706
rect 48446 -7764 48458 -7706
rect 49928 -7756 49940 -7664
rect 66588 -7756 66600 -7664
rect 49928 -7762 66600 -7756
rect 68108 -7710 68304 -7704
rect 48262 -7770 48458 -7764
rect 68108 -7768 68120 -7710
rect 68292 -7768 68304 -7710
rect 68914 -7756 68924 -6672
rect 69290 -7756 69300 -6672
rect 68108 -7774 68304 -7768
<< via1 >>
rect 47260 -6264 47620 -5190
rect 48286 -5236 48458 -5178
rect 49920 -5280 66568 -5188
rect 68070 -5236 68242 -5178
rect 50087 -5494 50139 -5442
rect 50277 -5493 50329 -5441
rect 50470 -5496 50522 -5444
rect 50662 -5491 50714 -5439
rect 50854 -5495 50906 -5443
rect 51046 -5490 51098 -5438
rect 51238 -5491 51290 -5439
rect 51428 -5490 51480 -5438
rect 51622 -5501 51674 -5449
rect 51811 -5499 51863 -5447
rect 52001 -5499 52053 -5447
rect 52200 -5500 52252 -5448
rect 52392 -5499 52444 -5447
rect 52582 -5500 52634 -5448
rect 52774 -5493 52826 -5441
rect 52966 -5495 53018 -5443
rect 53159 -5494 53211 -5442
rect 53351 -5492 53403 -5440
rect 53542 -5492 53594 -5440
rect 53736 -5497 53788 -5445
rect 53927 -5493 53979 -5441
rect 54119 -5489 54171 -5437
rect 54312 -5493 54364 -5441
rect 54504 -5493 54556 -5441
rect 54697 -5494 54749 -5442
rect 54889 -5492 54941 -5440
rect 55080 -5491 55132 -5439
rect 55271 -5490 55323 -5438
rect 55464 -5490 55516 -5438
rect 55655 -5499 55707 -5447
rect 55846 -5500 55898 -5448
rect 56036 -5501 56088 -5449
rect 56230 -5505 56282 -5453
rect 56422 -5507 56474 -5455
rect 56616 -5506 56668 -5454
rect 56808 -5503 56860 -5451
rect 56997 -5500 57049 -5448
rect 57191 -5498 57243 -5446
rect 57384 -5499 57436 -5447
rect 57577 -5500 57629 -5448
rect 57766 -5500 57818 -5448
rect 57959 -5500 58011 -5448
rect 58151 -5500 58203 -5448
rect 58342 -5500 58394 -5448
rect 58535 -5500 58587 -5448
rect 58726 -5499 58778 -5447
rect 58921 -5500 58973 -5448
rect 59110 -5500 59162 -5448
rect 59303 -5500 59355 -5448
rect 59495 -5500 59547 -5448
rect 59686 -5500 59738 -5448
rect 59878 -5500 59930 -5448
rect 60071 -5500 60123 -5448
rect 60260 -5501 60312 -5449
rect 60454 -5500 60506 -5448
rect 60645 -5500 60697 -5448
rect 60838 -5500 60890 -5448
rect 61030 -5500 61082 -5448
rect 61222 -5501 61274 -5449
rect 61415 -5499 61467 -5447
rect 61605 -5499 61657 -5447
rect 61798 -5501 61850 -5449
rect 61990 -5500 62042 -5448
rect 62183 -5499 62235 -5447
rect 62374 -5499 62426 -5447
rect 62566 -5500 62618 -5448
rect 62757 -5500 62809 -5448
rect 62949 -5500 63001 -5448
rect 63143 -5499 63195 -5447
rect 63335 -5500 63387 -5448
rect 63525 -5501 63577 -5449
rect 63716 -5502 63768 -5450
rect 63909 -5500 63961 -5448
rect 64102 -5499 64154 -5447
rect 64295 -5500 64347 -5448
rect 64486 -5500 64538 -5448
rect 64677 -5500 64729 -5448
rect 64870 -5500 64922 -5448
rect 65063 -5500 65115 -5448
rect 65254 -5500 65306 -5448
rect 65445 -5499 65497 -5447
rect 65636 -5499 65688 -5447
rect 65829 -5500 65881 -5448
rect 66023 -5500 66075 -5448
rect 66211 -5501 66263 -5449
rect 66405 -5509 66457 -5457
rect 49991 -5637 50043 -5585
rect 50182 -5639 50234 -5587
rect 50374 -5638 50426 -5586
rect 50566 -5641 50618 -5589
rect 50760 -5640 50812 -5588
rect 50950 -5640 51002 -5588
rect 51145 -5638 51197 -5586
rect 51336 -5637 51388 -5585
rect 51531 -5639 51583 -5587
rect 51721 -5639 51773 -5587
rect 51911 -5638 51963 -5586
rect 52104 -5637 52156 -5585
rect 52295 -5637 52347 -5585
rect 52491 -5639 52543 -5587
rect 52680 -5639 52732 -5587
rect 52874 -5639 52926 -5587
rect 53063 -5639 53115 -5587
rect 53255 -5640 53307 -5588
rect 53448 -5640 53500 -5588
rect 53639 -5640 53691 -5588
rect 53831 -5639 53883 -5587
rect 54023 -5640 54075 -5588
rect 54216 -5640 54268 -5588
rect 54407 -5640 54459 -5588
rect 54599 -5639 54651 -5587
rect 54792 -5640 54844 -5588
rect 54984 -5640 55036 -5588
rect 55175 -5640 55227 -5588
rect 55366 -5640 55418 -5588
rect 55558 -5640 55610 -5588
rect 55751 -5639 55803 -5587
rect 55942 -5639 55994 -5587
rect 56136 -5640 56188 -5588
rect 56328 -5640 56380 -5588
rect 56520 -5640 56572 -5588
rect 56712 -5640 56764 -5588
rect 56904 -5640 56956 -5588
rect 57096 -5640 57148 -5588
rect 57288 -5640 57340 -5588
rect 57479 -5640 57531 -5588
rect 57671 -5640 57723 -5588
rect 57864 -5640 57916 -5588
rect 58056 -5640 58108 -5588
rect 58248 -5640 58300 -5588
rect 58439 -5640 58491 -5588
rect 58631 -5640 58683 -5588
rect 58822 -5640 58874 -5588
rect 59013 -5640 59065 -5588
rect 59207 -5640 59259 -5588
rect 59399 -5640 59451 -5588
rect 59592 -5639 59644 -5587
rect 59783 -5640 59835 -5588
rect 59975 -5640 60027 -5588
rect 60168 -5640 60220 -5588
rect 60360 -5640 60412 -5588
rect 60553 -5639 60605 -5587
rect 60744 -5640 60796 -5588
rect 60936 -5640 60988 -5588
rect 61127 -5640 61179 -5588
rect 61319 -5640 61371 -5588
rect 61511 -5640 61563 -5588
rect 61704 -5640 61756 -5588
rect 61895 -5640 61947 -5588
rect 62087 -5640 62139 -5588
rect 62279 -5639 62331 -5587
rect 62471 -5640 62523 -5588
rect 62661 -5640 62713 -5588
rect 62855 -5640 62907 -5588
rect 63047 -5639 63099 -5587
rect 63238 -5640 63290 -5588
rect 63431 -5640 63483 -5588
rect 63622 -5639 63674 -5587
rect 63814 -5640 63866 -5588
rect 64005 -5640 64057 -5588
rect 64199 -5639 64251 -5587
rect 64390 -5640 64442 -5588
rect 64582 -5640 64634 -5588
rect 64774 -5640 64826 -5588
rect 64966 -5640 65018 -5588
rect 65159 -5640 65211 -5588
rect 65350 -5640 65402 -5588
rect 65543 -5639 65595 -5587
rect 65734 -5640 65786 -5588
rect 65927 -5640 65979 -5588
rect 66118 -5640 66170 -5588
rect 66309 -5638 66361 -5586
rect 66504 -5640 66556 -5588
rect 49430 -6126 49482 -6074
rect 51842 -6176 51898 -6120
rect 52047 -6123 52099 -6071
rect 52237 -6122 52289 -6070
rect 52429 -6121 52481 -6069
rect 52620 -6121 52672 -6069
rect 52814 -6121 52866 -6069
rect 53004 -6122 53056 -6070
rect 53198 -6121 53250 -6069
rect 53390 -6121 53442 -6069
rect 53581 -6122 53633 -6070
rect 53776 -6122 53828 -6070
rect 53966 -6122 54018 -6070
rect 54157 -6122 54209 -6070
rect 54349 -6122 54401 -6070
rect 54542 -6121 54594 -6069
rect 54734 -6122 54786 -6070
rect 54926 -6122 54978 -6070
rect 55119 -6122 55171 -6070
rect 55310 -6121 55362 -6069
rect 55502 -6122 55554 -6070
rect 55694 -6121 55746 -6069
rect 55886 -6121 55938 -6069
rect 56077 -6122 56129 -6070
rect 56270 -6121 56322 -6069
rect 56462 -6121 56514 -6069
rect 56656 -6122 56708 -6070
rect 56847 -6123 56899 -6071
rect 57036 -6122 57088 -6070
rect 57229 -6122 57281 -6070
rect 57422 -6122 57474 -6070
rect 57613 -6121 57665 -6069
rect 57804 -6121 57856 -6069
rect 58241 -6122 58293 -6070
rect 58431 -6121 58483 -6069
rect 58623 -6120 58675 -6068
rect 58814 -6120 58866 -6068
rect 59008 -6120 59060 -6068
rect 59198 -6121 59250 -6069
rect 59392 -6120 59444 -6068
rect 59584 -6120 59636 -6068
rect 59775 -6121 59827 -6069
rect 59970 -6121 60022 -6069
rect 60160 -6121 60212 -6069
rect 60351 -6121 60403 -6069
rect 60543 -6121 60595 -6069
rect 60736 -6120 60788 -6068
rect 60928 -6121 60980 -6069
rect 61120 -6121 61172 -6069
rect 61313 -6121 61365 -6069
rect 61504 -6120 61556 -6068
rect 61696 -6121 61748 -6069
rect 61888 -6120 61940 -6068
rect 62080 -6120 62132 -6068
rect 62271 -6121 62323 -6069
rect 62464 -6120 62516 -6068
rect 62656 -6120 62708 -6068
rect 62850 -6121 62902 -6069
rect 63041 -6122 63093 -6070
rect 63230 -6121 63282 -6069
rect 63423 -6121 63475 -6069
rect 63616 -6121 63668 -6069
rect 63807 -6120 63859 -6068
rect 63998 -6120 64050 -6068
rect 51942 -6262 51998 -6206
rect 52134 -6264 52190 -6208
rect 52328 -6266 52384 -6210
rect 52524 -6266 52580 -6210
rect 52714 -6270 52770 -6214
rect 52906 -6266 52962 -6210
rect 53100 -6268 53156 -6212
rect 53288 -6266 53344 -6210
rect 53480 -6268 53536 -6212
rect 53672 -6264 53728 -6208
rect 53870 -6266 53926 -6210
rect 54058 -6268 54114 -6212
rect 54252 -6266 54308 -6210
rect 54440 -6264 54496 -6208
rect 54632 -6270 54688 -6214
rect 54826 -6268 54882 -6212
rect 55016 -6268 55072 -6212
rect 55212 -6268 55268 -6212
rect 55402 -6268 55458 -6212
rect 55594 -6266 55650 -6210
rect 55786 -6264 55842 -6208
rect 55978 -6266 56034 -6210
rect 56172 -6264 56228 -6208
rect 56362 -6268 56418 -6212
rect 56558 -6266 56614 -6210
rect 56746 -6266 56802 -6210
rect 56940 -6266 56996 -6210
rect 57132 -6266 57188 -6210
rect 57318 -6270 57374 -6214
rect 57516 -6268 57572 -6212
rect 57702 -6268 57758 -6212
rect 58138 -6266 58194 -6210
rect 58330 -6268 58386 -6212
rect 58526 -6266 58582 -6210
rect 58714 -6268 58770 -6212
rect 58906 -6270 58962 -6214
rect 59100 -6268 59156 -6212
rect 59292 -6270 59348 -6214
rect 59484 -6268 59540 -6212
rect 59678 -6266 59734 -6210
rect 59868 -6266 59924 -6210
rect 60060 -6270 60116 -6214
rect 60252 -6270 60308 -6214
rect 60444 -6268 60500 -6212
rect 60638 -6268 60694 -6212
rect 60828 -6270 60884 -6214
rect 61018 -6268 61074 -6212
rect 61212 -6264 61268 -6208
rect 61404 -6270 61460 -6214
rect 61596 -6270 61652 -6214
rect 61786 -6270 61842 -6214
rect 61976 -6268 62032 -6212
rect 62174 -6266 62230 -6210
rect 62364 -6270 62420 -6214
rect 62554 -6268 62610 -6212
rect 62750 -6268 62806 -6212
rect 62938 -6266 62994 -6210
rect 63134 -6270 63190 -6214
rect 63322 -6268 63378 -6212
rect 63512 -6266 63568 -6210
rect 63710 -6268 63766 -6212
rect 63902 -6266 63958 -6210
rect 64128 -6232 64184 -6176
rect 51726 -6438 51782 -6382
rect 66918 -6002 66970 -5950
rect 68930 -6272 69296 -5188
rect 64236 -6456 64292 -6400
rect 47254 -7752 47614 -6678
rect 49436 -6924 49488 -6872
rect 52044 -6746 52100 -6690
rect 52238 -6746 52294 -6690
rect 52432 -6752 52488 -6696
rect 52622 -6748 52678 -6692
rect 52818 -6748 52874 -6692
rect 53006 -6748 53062 -6692
rect 53200 -6746 53256 -6690
rect 53394 -6746 53450 -6690
rect 53582 -6748 53638 -6692
rect 53774 -6746 53830 -6690
rect 53964 -6750 54020 -6694
rect 54156 -6748 54212 -6692
rect 54350 -6750 54406 -6694
rect 54542 -6746 54598 -6690
rect 54740 -6748 54796 -6692
rect 54926 -6746 54982 -6690
rect 55120 -6752 55176 -6696
rect 55310 -6748 55366 -6692
rect 55502 -6752 55558 -6696
rect 55690 -6746 55746 -6690
rect 55886 -6750 55942 -6694
rect 56078 -6744 56134 -6688
rect 56272 -6748 56328 -6692
rect 56460 -6750 56516 -6694
rect 56658 -6750 56714 -6694
rect 56848 -6746 56904 -6690
rect 57038 -6752 57094 -6696
rect 57228 -6746 57284 -6690
rect 57422 -6752 57478 -6696
rect 57608 -6748 57664 -6692
rect 57806 -6750 57862 -6694
rect 58230 -6750 58286 -6694
rect 58420 -6748 58476 -6692
rect 58612 -6754 58668 -6698
rect 58802 -6748 58858 -6692
rect 58996 -6750 59052 -6694
rect 59190 -6746 59246 -6690
rect 59382 -6750 59438 -6694
rect 59572 -6748 59628 -6692
rect 59764 -6750 59820 -6694
rect 59960 -6746 60016 -6690
rect 60154 -6748 60210 -6692
rect 60342 -6746 60398 -6690
rect 60534 -6752 60590 -6696
rect 60726 -6744 60782 -6688
rect 60918 -6750 60974 -6694
rect 61110 -6746 61166 -6690
rect 61300 -6750 61356 -6694
rect 61492 -6746 61548 -6690
rect 61688 -6752 61744 -6696
rect 61874 -6746 61930 -6690
rect 62070 -6748 62126 -6692
rect 62260 -6746 62316 -6690
rect 62456 -6748 62512 -6692
rect 62644 -6746 62700 -6690
rect 62840 -6746 62896 -6690
rect 63028 -6748 63084 -6692
rect 63220 -6748 63276 -6692
rect 63412 -6748 63468 -6692
rect 63608 -6746 63664 -6690
rect 63796 -6744 63852 -6688
rect 63992 -6746 64048 -6690
rect 51950 -6880 52002 -6828
rect 52142 -6880 52194 -6828
rect 52335 -6880 52387 -6828
rect 52527 -6880 52579 -6828
rect 52720 -6880 52772 -6828
rect 52912 -6879 52964 -6827
rect 53103 -6880 53155 -6828
rect 53295 -6880 53347 -6828
rect 53487 -6879 53539 -6827
rect 53679 -6879 53731 -6827
rect 53871 -6880 53923 -6828
rect 54063 -6879 54115 -6827
rect 54255 -6880 54307 -6828
rect 54446 -6879 54498 -6827
rect 54640 -6880 54692 -6828
rect 54830 -6880 54882 -6828
rect 55022 -6880 55074 -6828
rect 55215 -6880 55267 -6828
rect 55406 -6880 55458 -6828
rect 55599 -6879 55651 -6827
rect 55792 -6880 55844 -6828
rect 55983 -6880 56035 -6828
rect 56176 -6880 56228 -6828
rect 56366 -6880 56418 -6828
rect 56560 -6879 56612 -6827
rect 56749 -6880 56801 -6828
rect 56942 -6880 56994 -6828
rect 57135 -6880 57187 -6828
rect 57325 -6880 57377 -6828
rect 57518 -6879 57570 -6827
rect 57707 -6879 57759 -6827
rect 58138 -6879 58190 -6827
rect 58330 -6879 58382 -6827
rect 58523 -6879 58575 -6827
rect 58715 -6879 58767 -6827
rect 58908 -6879 58960 -6827
rect 59100 -6878 59152 -6826
rect 59291 -6879 59343 -6827
rect 59483 -6879 59535 -6827
rect 59675 -6878 59727 -6826
rect 59867 -6878 59919 -6826
rect 60059 -6879 60111 -6827
rect 60251 -6878 60303 -6826
rect 60443 -6879 60495 -6827
rect 60634 -6878 60686 -6826
rect 60828 -6879 60880 -6827
rect 61018 -6879 61070 -6827
rect 61210 -6879 61262 -6827
rect 61403 -6879 61455 -6827
rect 61594 -6879 61646 -6827
rect 61787 -6878 61839 -6826
rect 61980 -6879 62032 -6827
rect 62171 -6879 62223 -6827
rect 62364 -6879 62416 -6827
rect 62554 -6879 62606 -6827
rect 62748 -6878 62800 -6826
rect 62937 -6879 62989 -6827
rect 63130 -6879 63182 -6827
rect 63323 -6879 63375 -6827
rect 63513 -6879 63565 -6827
rect 63706 -6878 63758 -6826
rect 63895 -6878 63947 -6826
rect 66912 -6902 66964 -6850
rect 50087 -7354 50139 -7302
rect 50277 -7353 50329 -7301
rect 50470 -7356 50522 -7304
rect 50662 -7351 50714 -7299
rect 50854 -7355 50906 -7303
rect 51046 -7350 51098 -7298
rect 51238 -7351 51290 -7299
rect 51428 -7350 51480 -7298
rect 51622 -7361 51674 -7309
rect 51811 -7359 51863 -7307
rect 52001 -7359 52053 -7307
rect 52200 -7360 52252 -7308
rect 52392 -7359 52444 -7307
rect 52582 -7360 52634 -7308
rect 52774 -7353 52826 -7301
rect 52966 -7355 53018 -7303
rect 53159 -7354 53211 -7302
rect 53351 -7352 53403 -7300
rect 53542 -7352 53594 -7300
rect 53736 -7357 53788 -7305
rect 53927 -7353 53979 -7301
rect 54119 -7349 54171 -7297
rect 54312 -7353 54364 -7301
rect 54504 -7353 54556 -7301
rect 54697 -7354 54749 -7302
rect 54889 -7352 54941 -7300
rect 55080 -7351 55132 -7299
rect 55271 -7350 55323 -7298
rect 55464 -7350 55516 -7298
rect 55655 -7359 55707 -7307
rect 55846 -7360 55898 -7308
rect 56036 -7361 56088 -7309
rect 56230 -7365 56282 -7313
rect 56422 -7367 56474 -7315
rect 56616 -7366 56668 -7314
rect 56808 -7363 56860 -7311
rect 56997 -7360 57049 -7308
rect 57191 -7358 57243 -7306
rect 57384 -7359 57436 -7307
rect 57577 -7360 57629 -7308
rect 57766 -7360 57818 -7308
rect 57959 -7360 58011 -7308
rect 58151 -7360 58203 -7308
rect 58342 -7360 58394 -7308
rect 58535 -7360 58587 -7308
rect 58726 -7359 58778 -7307
rect 58921 -7360 58973 -7308
rect 59110 -7360 59162 -7308
rect 59303 -7360 59355 -7308
rect 59495 -7360 59547 -7308
rect 59686 -7360 59738 -7308
rect 59878 -7360 59930 -7308
rect 60071 -7360 60123 -7308
rect 60260 -7361 60312 -7309
rect 60454 -7360 60506 -7308
rect 60645 -7360 60697 -7308
rect 60838 -7360 60890 -7308
rect 61030 -7360 61082 -7308
rect 61222 -7361 61274 -7309
rect 61415 -7359 61467 -7307
rect 61605 -7359 61657 -7307
rect 61798 -7361 61850 -7309
rect 61990 -7360 62042 -7308
rect 62183 -7359 62235 -7307
rect 62374 -7359 62426 -7307
rect 62566 -7360 62618 -7308
rect 62757 -7360 62809 -7308
rect 62949 -7360 63001 -7308
rect 63143 -7359 63195 -7307
rect 63335 -7360 63387 -7308
rect 63525 -7361 63577 -7309
rect 63716 -7362 63768 -7310
rect 63909 -7360 63961 -7308
rect 64102 -7359 64154 -7307
rect 64295 -7360 64347 -7308
rect 64486 -7360 64538 -7308
rect 64677 -7360 64729 -7308
rect 64870 -7360 64922 -7308
rect 65063 -7360 65115 -7308
rect 65254 -7360 65306 -7308
rect 65445 -7359 65497 -7307
rect 65636 -7359 65688 -7307
rect 65829 -7360 65881 -7308
rect 66023 -7360 66075 -7308
rect 66211 -7361 66263 -7309
rect 66405 -7369 66457 -7317
rect 49991 -7497 50043 -7445
rect 50182 -7499 50234 -7447
rect 50374 -7498 50426 -7446
rect 50566 -7501 50618 -7449
rect 50760 -7500 50812 -7448
rect 50950 -7500 51002 -7448
rect 51145 -7498 51197 -7446
rect 51336 -7497 51388 -7445
rect 51531 -7499 51583 -7447
rect 51721 -7499 51773 -7447
rect 51911 -7498 51963 -7446
rect 52104 -7497 52156 -7445
rect 52295 -7497 52347 -7445
rect 52491 -7499 52543 -7447
rect 52680 -7499 52732 -7447
rect 52874 -7499 52926 -7447
rect 53063 -7499 53115 -7447
rect 53255 -7500 53307 -7448
rect 53448 -7500 53500 -7448
rect 53639 -7500 53691 -7448
rect 53831 -7499 53883 -7447
rect 54023 -7500 54075 -7448
rect 54216 -7500 54268 -7448
rect 54407 -7500 54459 -7448
rect 54599 -7499 54651 -7447
rect 54792 -7500 54844 -7448
rect 54984 -7500 55036 -7448
rect 55175 -7500 55227 -7448
rect 55366 -7500 55418 -7448
rect 55558 -7500 55610 -7448
rect 55751 -7499 55803 -7447
rect 55942 -7499 55994 -7447
rect 56136 -7500 56188 -7448
rect 56328 -7500 56380 -7448
rect 56520 -7500 56572 -7448
rect 56712 -7500 56764 -7448
rect 56904 -7500 56956 -7448
rect 57096 -7500 57148 -7448
rect 57288 -7500 57340 -7448
rect 57479 -7500 57531 -7448
rect 57671 -7500 57723 -7448
rect 57864 -7500 57916 -7448
rect 58056 -7500 58108 -7448
rect 58248 -7500 58300 -7448
rect 58439 -7500 58491 -7448
rect 58631 -7500 58683 -7448
rect 58822 -7500 58874 -7448
rect 59013 -7500 59065 -7448
rect 59207 -7500 59259 -7448
rect 59399 -7500 59451 -7448
rect 59592 -7499 59644 -7447
rect 59783 -7500 59835 -7448
rect 59975 -7500 60027 -7448
rect 60168 -7500 60220 -7448
rect 60360 -7500 60412 -7448
rect 60553 -7499 60605 -7447
rect 60744 -7500 60796 -7448
rect 60936 -7500 60988 -7448
rect 61127 -7500 61179 -7448
rect 61319 -7500 61371 -7448
rect 61511 -7500 61563 -7448
rect 61704 -7500 61756 -7448
rect 61895 -7500 61947 -7448
rect 62087 -7500 62139 -7448
rect 62279 -7499 62331 -7447
rect 62471 -7500 62523 -7448
rect 62661 -7500 62713 -7448
rect 62855 -7500 62907 -7448
rect 63047 -7499 63099 -7447
rect 63238 -7500 63290 -7448
rect 63431 -7500 63483 -7448
rect 63622 -7499 63674 -7447
rect 63814 -7500 63866 -7448
rect 64005 -7500 64057 -7448
rect 64199 -7499 64251 -7447
rect 64390 -7500 64442 -7448
rect 64582 -7500 64634 -7448
rect 64774 -7500 64826 -7448
rect 64966 -7500 65018 -7448
rect 65159 -7500 65211 -7448
rect 65350 -7500 65402 -7448
rect 65543 -7499 65595 -7447
rect 65734 -7500 65786 -7448
rect 65927 -7500 65979 -7448
rect 66118 -7500 66170 -7448
rect 66309 -7498 66361 -7446
rect 66504 -7500 66556 -7448
rect 48274 -7764 48446 -7706
rect 49940 -7756 66588 -7664
rect 68120 -7768 68292 -7710
rect 68924 -7756 69290 -6672
<< metal2 >>
rect 68894 -4738 69326 -4736
rect 68674 -4740 69326 -4738
rect 47224 -5130 69326 -4740
rect 47224 -5190 47652 -5130
rect 47224 -6264 47260 -5190
rect 47620 -6264 47652 -5190
rect 48286 -5178 48458 -5168
rect 68070 -5178 68242 -5168
rect 48286 -5246 48458 -5236
rect 49920 -5188 66568 -5178
rect 68070 -5246 68242 -5236
rect 68894 -5188 69326 -5130
rect 49920 -5290 66568 -5280
rect 50090 -5432 50160 -5290
rect 50087 -5440 50160 -5432
rect 50277 -5440 50329 -5431
rect 50470 -5440 50522 -5434
rect 50662 -5439 50714 -5430
rect 50087 -5441 50662 -5440
rect 50087 -5442 50277 -5441
rect 50139 -5470 50277 -5442
rect 50087 -5504 50139 -5494
rect 50329 -5444 50662 -5441
rect 50329 -5470 50470 -5444
rect 50277 -5503 50329 -5493
rect 50522 -5470 50662 -5444
rect 50470 -5506 50522 -5496
rect 50854 -5440 50906 -5433
rect 51046 -5438 51098 -5430
rect 50714 -5443 51046 -5440
rect 50714 -5470 50854 -5443
rect 50662 -5501 50714 -5491
rect 50906 -5470 51046 -5443
rect 50854 -5505 50906 -5495
rect 51238 -5439 51290 -5430
rect 51098 -5470 51238 -5440
rect 51046 -5500 51098 -5490
rect 51428 -5438 51480 -5430
rect 51290 -5470 51428 -5440
rect 51238 -5501 51290 -5491
rect 51622 -5440 51674 -5439
rect 51811 -5440 51863 -5437
rect 52001 -5440 52053 -5437
rect 52200 -5440 52252 -5438
rect 52392 -5440 52444 -5437
rect 52582 -5440 52634 -5438
rect 52774 -5440 52826 -5431
rect 52966 -5440 53018 -5433
rect 53159 -5440 53211 -5432
rect 53351 -5440 53403 -5430
rect 53542 -5440 53594 -5430
rect 53736 -5440 53788 -5435
rect 53927 -5440 53979 -5431
rect 54119 -5437 54171 -5430
rect 51480 -5441 53351 -5440
rect 51480 -5447 52774 -5441
rect 51480 -5449 51811 -5447
rect 51480 -5470 51622 -5449
rect 51428 -5500 51480 -5490
rect 51674 -5470 51811 -5449
rect 51622 -5511 51674 -5501
rect 51863 -5470 52001 -5447
rect 51811 -5509 51863 -5499
rect 52053 -5448 52392 -5447
rect 52053 -5470 52200 -5448
rect 52001 -5509 52053 -5499
rect 52252 -5470 52392 -5448
rect 52200 -5510 52252 -5500
rect 52444 -5448 52774 -5447
rect 52444 -5470 52582 -5448
rect 52392 -5509 52444 -5499
rect 52634 -5470 52774 -5448
rect 52582 -5510 52634 -5500
rect 52826 -5442 53351 -5441
rect 52826 -5443 53159 -5442
rect 52826 -5470 52966 -5443
rect 52774 -5503 52826 -5493
rect 53018 -5470 53159 -5443
rect 52966 -5505 53018 -5495
rect 53211 -5470 53351 -5442
rect 53159 -5504 53211 -5494
rect 53403 -5470 53542 -5440
rect 53351 -5502 53403 -5492
rect 53594 -5441 54119 -5440
rect 53594 -5445 53927 -5441
rect 53594 -5470 53736 -5445
rect 53542 -5502 53594 -5492
rect 53788 -5470 53927 -5445
rect 53736 -5507 53788 -5497
rect 53979 -5470 54119 -5441
rect 53927 -5503 53979 -5493
rect 54312 -5440 54364 -5431
rect 54504 -5440 54556 -5431
rect 54697 -5440 54749 -5432
rect 54889 -5440 54941 -5430
rect 55080 -5439 55132 -5430
rect 54171 -5441 54889 -5440
rect 54171 -5470 54312 -5441
rect 54119 -5499 54171 -5489
rect 54364 -5470 54504 -5441
rect 54312 -5503 54364 -5493
rect 54556 -5442 54889 -5441
rect 54556 -5470 54697 -5442
rect 54504 -5503 54556 -5493
rect 54749 -5470 54889 -5442
rect 54697 -5504 54749 -5494
rect 54941 -5470 55080 -5440
rect 54889 -5502 54941 -5492
rect 55271 -5438 55323 -5430
rect 55132 -5470 55271 -5440
rect 55080 -5501 55132 -5491
rect 55464 -5438 55516 -5430
rect 55323 -5470 55464 -5440
rect 55271 -5500 55323 -5490
rect 55655 -5440 55707 -5437
rect 55846 -5440 55898 -5438
rect 56036 -5440 56088 -5439
rect 56997 -5440 57049 -5438
rect 57191 -5440 57243 -5436
rect 57384 -5440 57436 -5437
rect 57577 -5440 57629 -5438
rect 57766 -5440 57818 -5438
rect 57959 -5440 58011 -5438
rect 58151 -5440 58203 -5438
rect 58342 -5440 58394 -5438
rect 58535 -5440 58587 -5438
rect 58726 -5440 58778 -5437
rect 58921 -5440 58973 -5438
rect 59110 -5440 59162 -5438
rect 59303 -5440 59355 -5438
rect 59495 -5440 59547 -5438
rect 59686 -5440 59738 -5438
rect 59878 -5440 59930 -5438
rect 60071 -5440 60123 -5438
rect 60260 -5440 60312 -5439
rect 60454 -5440 60506 -5438
rect 60645 -5440 60697 -5438
rect 60838 -5440 60890 -5438
rect 61030 -5440 61082 -5438
rect 61222 -5440 61274 -5439
rect 61415 -5440 61467 -5437
rect 61605 -5440 61657 -5437
rect 61798 -5440 61850 -5439
rect 61990 -5440 62042 -5438
rect 62183 -5440 62235 -5437
rect 62374 -5440 62426 -5437
rect 62566 -5440 62618 -5438
rect 62757 -5440 62809 -5438
rect 62949 -5440 63001 -5438
rect 63143 -5440 63195 -5437
rect 63335 -5440 63387 -5438
rect 63525 -5440 63577 -5439
rect 63909 -5440 63961 -5438
rect 64102 -5440 64154 -5437
rect 64295 -5440 64347 -5438
rect 64486 -5440 64538 -5438
rect 64677 -5440 64729 -5438
rect 64870 -5440 64922 -5438
rect 65063 -5440 65115 -5438
rect 65254 -5440 65306 -5438
rect 65445 -5440 65497 -5437
rect 65636 -5440 65688 -5437
rect 65829 -5440 65881 -5438
rect 66023 -5440 66075 -5438
rect 66211 -5440 66263 -5439
rect 66400 -5440 66470 -5290
rect 55516 -5446 66470 -5440
rect 55516 -5447 57191 -5446
rect 55516 -5470 55655 -5447
rect 55464 -5500 55516 -5490
rect 55707 -5448 57191 -5447
rect 55707 -5470 55846 -5448
rect 55655 -5509 55707 -5499
rect 55898 -5449 56997 -5448
rect 55898 -5470 56036 -5449
rect 55846 -5510 55898 -5500
rect 56088 -5451 56997 -5449
rect 56088 -5453 56808 -5451
rect 56088 -5470 56230 -5453
rect 56036 -5511 56088 -5501
rect 56282 -5454 56808 -5453
rect 56282 -5455 56616 -5454
rect 56282 -5470 56422 -5455
rect 56230 -5515 56282 -5505
rect 56474 -5470 56616 -5455
rect 56422 -5517 56474 -5507
rect 56668 -5470 56808 -5454
rect 56616 -5516 56668 -5506
rect 56860 -5470 56997 -5451
rect 56808 -5513 56860 -5503
rect 57049 -5470 57191 -5448
rect 56997 -5510 57049 -5500
rect 57243 -5447 66470 -5446
rect 57243 -5470 57384 -5447
rect 57191 -5508 57243 -5498
rect 57436 -5448 58726 -5447
rect 57436 -5470 57577 -5448
rect 57384 -5509 57436 -5499
rect 57629 -5470 57766 -5448
rect 57577 -5510 57629 -5500
rect 57818 -5470 57959 -5448
rect 57766 -5510 57818 -5500
rect 58011 -5470 58151 -5448
rect 57959 -5510 58011 -5500
rect 58203 -5470 58342 -5448
rect 58151 -5510 58203 -5500
rect 58394 -5470 58535 -5448
rect 58342 -5510 58394 -5500
rect 58587 -5470 58726 -5448
rect 58535 -5510 58587 -5500
rect 58778 -5448 61415 -5447
rect 58778 -5470 58921 -5448
rect 58726 -5509 58778 -5499
rect 58973 -5470 59110 -5448
rect 58921 -5510 58973 -5500
rect 59162 -5470 59303 -5448
rect 59110 -5510 59162 -5500
rect 59355 -5470 59495 -5448
rect 59303 -5510 59355 -5500
rect 59547 -5470 59686 -5448
rect 59495 -5510 59547 -5500
rect 59738 -5470 59878 -5448
rect 59686 -5510 59738 -5500
rect 59930 -5470 60071 -5448
rect 59878 -5510 59930 -5500
rect 60123 -5449 60454 -5448
rect 60123 -5470 60260 -5449
rect 60071 -5510 60123 -5500
rect 60312 -5470 60454 -5449
rect 60260 -5511 60312 -5501
rect 60506 -5470 60645 -5448
rect 60454 -5510 60506 -5500
rect 60697 -5470 60838 -5448
rect 60645 -5510 60697 -5500
rect 60890 -5470 61030 -5448
rect 60838 -5510 60890 -5500
rect 61082 -5449 61415 -5448
rect 61082 -5470 61222 -5449
rect 61030 -5510 61082 -5500
rect 61274 -5470 61415 -5449
rect 61222 -5511 61274 -5501
rect 61467 -5470 61605 -5447
rect 61415 -5509 61467 -5499
rect 61657 -5448 62183 -5447
rect 61657 -5449 61990 -5448
rect 61657 -5470 61798 -5449
rect 61605 -5509 61657 -5499
rect 61850 -5470 61990 -5449
rect 61798 -5511 61850 -5501
rect 62042 -5470 62183 -5448
rect 61990 -5510 62042 -5500
rect 62235 -5470 62374 -5447
rect 62183 -5509 62235 -5499
rect 62426 -5448 63143 -5447
rect 62426 -5470 62566 -5448
rect 62374 -5509 62426 -5499
rect 62618 -5470 62757 -5448
rect 62566 -5510 62618 -5500
rect 62809 -5470 62949 -5448
rect 62757 -5510 62809 -5500
rect 63001 -5470 63143 -5448
rect 62949 -5510 63001 -5500
rect 63195 -5448 64102 -5447
rect 63195 -5470 63335 -5448
rect 63143 -5509 63195 -5499
rect 63387 -5449 63909 -5448
rect 63387 -5470 63525 -5449
rect 63335 -5510 63387 -5500
rect 63577 -5450 63909 -5449
rect 63577 -5470 63716 -5450
rect 63525 -5511 63577 -5501
rect 63768 -5470 63909 -5450
rect 63716 -5512 63768 -5502
rect 63961 -5470 64102 -5448
rect 63909 -5510 63961 -5500
rect 64154 -5448 65445 -5447
rect 64154 -5470 64295 -5448
rect 64102 -5509 64154 -5499
rect 64347 -5470 64486 -5448
rect 64295 -5510 64347 -5500
rect 64538 -5470 64677 -5448
rect 64486 -5510 64538 -5500
rect 64729 -5470 64870 -5448
rect 64677 -5510 64729 -5500
rect 64922 -5470 65063 -5448
rect 64870 -5510 64922 -5500
rect 65115 -5470 65254 -5448
rect 65063 -5510 65115 -5500
rect 65306 -5470 65445 -5448
rect 65254 -5510 65306 -5500
rect 65497 -5470 65636 -5447
rect 65445 -5509 65497 -5499
rect 65688 -5448 66470 -5447
rect 65688 -5470 65829 -5448
rect 65636 -5509 65688 -5499
rect 65881 -5470 66023 -5448
rect 65829 -5510 65881 -5500
rect 66075 -5449 66470 -5448
rect 66075 -5470 66211 -5449
rect 66023 -5510 66075 -5500
rect 66263 -5457 66470 -5449
rect 66263 -5470 66405 -5457
rect 66211 -5511 66263 -5501
rect 66457 -5470 66470 -5457
rect 66405 -5519 66457 -5509
rect 49991 -5585 50043 -5575
rect 50182 -5587 50234 -5577
rect 50043 -5630 50182 -5600
rect 49991 -5647 50043 -5637
rect 50374 -5586 50426 -5576
rect 50234 -5630 50374 -5600
rect 50182 -5649 50234 -5639
rect 50566 -5589 50618 -5579
rect 50426 -5630 50566 -5600
rect 50374 -5648 50426 -5638
rect 50760 -5588 50812 -5578
rect 50618 -5630 50760 -5600
rect 50566 -5651 50618 -5641
rect 50950 -5588 51002 -5578
rect 50812 -5630 50950 -5600
rect 50760 -5650 50812 -5640
rect 51145 -5586 51197 -5576
rect 51002 -5630 51145 -5600
rect 50950 -5650 51002 -5640
rect 51336 -5585 51388 -5575
rect 51197 -5630 51336 -5600
rect 51145 -5648 51197 -5638
rect 51531 -5587 51583 -5577
rect 51388 -5630 51531 -5600
rect 51336 -5647 51388 -5637
rect 51721 -5587 51773 -5577
rect 51583 -5630 51721 -5600
rect 51531 -5649 51583 -5639
rect 51911 -5586 51963 -5576
rect 51773 -5630 51911 -5600
rect 51721 -5649 51773 -5639
rect 52104 -5585 52156 -5575
rect 51963 -5630 52104 -5600
rect 51911 -5648 51963 -5638
rect 52050 -5637 52104 -5630
rect 52295 -5585 52347 -5575
rect 52156 -5630 52295 -5600
rect 52050 -5647 52156 -5637
rect 52491 -5587 52543 -5577
rect 52347 -5630 52491 -5600
rect 52295 -5647 52347 -5637
rect 52430 -5639 52491 -5630
rect 52680 -5587 52732 -5577
rect 52543 -5630 52680 -5600
rect 52050 -5966 52110 -5647
rect 52430 -5649 52543 -5639
rect 52874 -5587 52926 -5577
rect 52732 -5630 52874 -5600
rect 52680 -5649 52732 -5639
rect 52820 -5639 52874 -5630
rect 53063 -5587 53115 -5577
rect 52926 -5630 53063 -5600
rect 52820 -5649 52926 -5639
rect 53255 -5588 53307 -5578
rect 53115 -5630 53255 -5600
rect 53063 -5649 53115 -5639
rect 53200 -5640 53255 -5630
rect 53448 -5588 53500 -5578
rect 53307 -5630 53448 -5600
rect 52430 -5966 52490 -5649
rect 52820 -5966 52880 -5649
rect 53200 -5650 53307 -5640
rect 53639 -5588 53691 -5578
rect 53500 -5630 53639 -5600
rect 53448 -5650 53500 -5640
rect 53580 -5640 53639 -5630
rect 53831 -5587 53883 -5577
rect 53691 -5630 53831 -5600
rect 53580 -5650 53691 -5640
rect 54023 -5588 54075 -5578
rect 53883 -5630 54023 -5600
rect 53831 -5649 53883 -5639
rect 53970 -5640 54023 -5630
rect 54216 -5588 54268 -5578
rect 54075 -5630 54216 -5600
rect 53970 -5650 54075 -5640
rect 54407 -5588 54459 -5578
rect 54268 -5630 54407 -5600
rect 54216 -5650 54268 -5640
rect 54350 -5640 54407 -5630
rect 54599 -5587 54651 -5577
rect 54459 -5630 54599 -5600
rect 54350 -5650 54459 -5640
rect 54792 -5588 54844 -5578
rect 54651 -5630 54792 -5600
rect 54599 -5649 54651 -5639
rect 54740 -5640 54792 -5630
rect 54984 -5588 55036 -5578
rect 54844 -5630 54984 -5600
rect 54740 -5650 54844 -5640
rect 55175 -5588 55227 -5578
rect 55036 -5630 55175 -5600
rect 54984 -5650 55036 -5640
rect 55120 -5640 55175 -5630
rect 55366 -5588 55418 -5578
rect 55227 -5630 55366 -5600
rect 55120 -5650 55227 -5640
rect 55558 -5588 55610 -5578
rect 55418 -5630 55558 -5600
rect 55366 -5650 55418 -5640
rect 55500 -5640 55558 -5630
rect 55751 -5587 55803 -5577
rect 55610 -5630 55751 -5600
rect 55500 -5650 55610 -5640
rect 55942 -5587 55994 -5577
rect 55803 -5630 55942 -5600
rect 55751 -5649 55803 -5639
rect 55890 -5639 55942 -5630
rect 56136 -5588 56188 -5578
rect 55994 -5630 56136 -5600
rect 55890 -5649 55994 -5639
rect 56328 -5588 56380 -5578
rect 56188 -5630 56328 -5600
rect 53200 -5966 53260 -5650
rect 53580 -5966 53640 -5650
rect 53970 -5966 54030 -5650
rect 54350 -5966 54410 -5650
rect 54740 -5966 54800 -5650
rect 55120 -5966 55180 -5650
rect 55500 -5966 55560 -5650
rect 55890 -5966 55950 -5649
rect 56136 -5650 56188 -5640
rect 56270 -5640 56328 -5630
rect 56520 -5588 56572 -5578
rect 56380 -5630 56520 -5600
rect 56270 -5650 56380 -5640
rect 56712 -5588 56764 -5578
rect 56572 -5630 56712 -5600
rect 56520 -5650 56572 -5640
rect 56660 -5640 56712 -5630
rect 56904 -5588 56956 -5578
rect 56764 -5630 56904 -5600
rect 56660 -5650 56764 -5640
rect 57096 -5588 57148 -5578
rect 56956 -5630 57096 -5600
rect 56904 -5650 56956 -5640
rect 57040 -5640 57096 -5630
rect 57288 -5588 57340 -5578
rect 57148 -5630 57288 -5600
rect 57040 -5650 57148 -5640
rect 57479 -5588 57531 -5578
rect 57340 -5630 57479 -5600
rect 57288 -5650 57340 -5640
rect 57420 -5640 57479 -5630
rect 57671 -5588 57723 -5578
rect 57531 -5630 57671 -5600
rect 57420 -5650 57531 -5640
rect 57864 -5588 57916 -5578
rect 57723 -5630 57864 -5600
rect 57671 -5650 57723 -5640
rect 57810 -5640 57864 -5630
rect 58056 -5588 58108 -5578
rect 57916 -5630 58056 -5600
rect 57810 -5650 57916 -5640
rect 58248 -5588 58300 -5578
rect 58108 -5630 58248 -5600
rect 58056 -5650 58108 -5640
rect 58240 -5640 58248 -5630
rect 58439 -5588 58491 -5578
rect 58300 -5630 58439 -5600
rect 56270 -5966 56330 -5650
rect 56660 -5966 56720 -5650
rect 57040 -5966 57100 -5650
rect 57420 -5966 57480 -5650
rect 57810 -5966 57870 -5650
rect 58240 -5966 58300 -5640
rect 58631 -5588 58683 -5578
rect 58491 -5630 58631 -5600
rect 58439 -5650 58491 -5640
rect 58620 -5640 58631 -5630
rect 58822 -5588 58874 -5578
rect 58683 -5630 58822 -5600
rect 58620 -5650 58683 -5640
rect 59013 -5588 59065 -5578
rect 58874 -5630 59013 -5600
rect 58822 -5650 58874 -5640
rect 59010 -5640 59013 -5630
rect 59207 -5588 59259 -5578
rect 59065 -5630 59207 -5600
rect 59065 -5640 59070 -5630
rect 58620 -5966 58680 -5650
rect 59010 -5966 59070 -5640
rect 59399 -5588 59451 -5578
rect 59259 -5630 59399 -5600
rect 59207 -5650 59259 -5640
rect 59592 -5587 59644 -5577
rect 59451 -5630 59592 -5600
rect 59451 -5640 59460 -5630
rect 59399 -5650 59460 -5640
rect 59783 -5588 59835 -5578
rect 59644 -5630 59783 -5600
rect 59592 -5649 59644 -5639
rect 59780 -5640 59783 -5630
rect 59975 -5588 60027 -5578
rect 59835 -5630 59975 -5600
rect 59835 -5640 59840 -5630
rect 59400 -5966 59460 -5650
rect 59780 -5966 59840 -5640
rect 60168 -5588 60220 -5578
rect 60027 -5630 60168 -5600
rect 59975 -5650 60027 -5640
rect 60160 -5640 60168 -5630
rect 60360 -5588 60412 -5578
rect 60220 -5630 60360 -5600
rect 60160 -5966 60220 -5640
rect 60553 -5587 60605 -5577
rect 60412 -5630 60553 -5600
rect 60360 -5650 60412 -5640
rect 60540 -5639 60553 -5630
rect 60744 -5588 60796 -5578
rect 60605 -5630 60744 -5600
rect 60540 -5649 60605 -5639
rect 60936 -5588 60988 -5578
rect 60796 -5630 60936 -5600
rect 60540 -5966 60600 -5649
rect 60744 -5650 60796 -5640
rect 60930 -5640 60936 -5630
rect 61127 -5588 61179 -5578
rect 60988 -5630 61127 -5600
rect 60988 -5640 60990 -5630
rect 60930 -5966 60990 -5640
rect 61319 -5588 61371 -5578
rect 61179 -5630 61319 -5600
rect 61127 -5650 61179 -5640
rect 61511 -5588 61563 -5578
rect 61371 -5630 61511 -5600
rect 61371 -5640 61380 -5630
rect 61319 -5650 61380 -5640
rect 61704 -5588 61756 -5578
rect 61563 -5630 61704 -5600
rect 61511 -5650 61563 -5640
rect 61700 -5640 61704 -5630
rect 61895 -5588 61947 -5578
rect 61756 -5630 61895 -5600
rect 61756 -5640 61760 -5630
rect 61320 -5966 61380 -5650
rect 61700 -5966 61760 -5640
rect 62087 -5588 62139 -5578
rect 61947 -5630 62087 -5600
rect 61895 -5650 61947 -5640
rect 62080 -5640 62087 -5630
rect 62279 -5587 62331 -5577
rect 62139 -5630 62279 -5600
rect 62139 -5640 62140 -5630
rect 62080 -5966 62140 -5640
rect 62471 -5588 62523 -5578
rect 62331 -5630 62471 -5600
rect 62279 -5649 62331 -5639
rect 62470 -5640 62471 -5630
rect 62661 -5588 62713 -5578
rect 62523 -5630 62661 -5600
rect 62523 -5640 62530 -5630
rect 62470 -5966 62530 -5640
rect 62855 -5588 62907 -5578
rect 62713 -5630 62855 -5600
rect 62661 -5650 62713 -5640
rect 62850 -5640 62855 -5630
rect 63047 -5587 63099 -5577
rect 62907 -5630 63047 -5600
rect 62907 -5640 62910 -5630
rect 62850 -5966 62910 -5640
rect 63238 -5588 63290 -5578
rect 63099 -5630 63238 -5600
rect 63047 -5649 63099 -5639
rect 63230 -5640 63238 -5630
rect 63431 -5588 63483 -5578
rect 63290 -5630 63431 -5600
rect 63230 -5966 63290 -5640
rect 63622 -5587 63674 -5577
rect 63483 -5630 63622 -5600
rect 63431 -5650 63483 -5640
rect 63620 -5639 63622 -5630
rect 63814 -5588 63866 -5578
rect 63674 -5630 63814 -5600
rect 63674 -5639 63680 -5630
rect 63620 -5966 63680 -5639
rect 64005 -5588 64057 -5578
rect 63866 -5630 64005 -5600
rect 63814 -5650 63866 -5640
rect 64000 -5640 64005 -5630
rect 64199 -5587 64251 -5577
rect 64057 -5630 64199 -5600
rect 64057 -5640 64060 -5630
rect 64000 -5966 64060 -5640
rect 64390 -5588 64442 -5578
rect 64251 -5630 64390 -5600
rect 64199 -5649 64251 -5639
rect 64582 -5588 64634 -5578
rect 64442 -5630 64582 -5600
rect 64390 -5650 64442 -5640
rect 64774 -5588 64826 -5578
rect 64634 -5630 64774 -5600
rect 64582 -5650 64634 -5640
rect 64966 -5588 65018 -5578
rect 64826 -5630 64966 -5600
rect 64774 -5650 64826 -5640
rect 65159 -5588 65211 -5578
rect 65018 -5630 65159 -5600
rect 64966 -5650 65018 -5640
rect 65350 -5588 65402 -5578
rect 65211 -5630 65350 -5600
rect 65159 -5650 65211 -5640
rect 65543 -5587 65595 -5577
rect 65402 -5630 65543 -5600
rect 65350 -5650 65402 -5640
rect 65734 -5588 65786 -5578
rect 65595 -5630 65734 -5600
rect 65543 -5649 65595 -5639
rect 65927 -5588 65979 -5578
rect 65786 -5630 65927 -5600
rect 65734 -5650 65786 -5640
rect 66118 -5588 66170 -5578
rect 65979 -5630 66118 -5600
rect 65927 -5650 65979 -5640
rect 66309 -5586 66361 -5576
rect 66170 -5630 66309 -5600
rect 66118 -5650 66170 -5640
rect 66504 -5588 66556 -5578
rect 66361 -5630 66504 -5600
rect 66309 -5648 66361 -5638
rect 66504 -5650 66556 -5640
rect 66918 -5950 66970 -5940
rect 52044 -6026 64072 -5966
rect 66918 -6012 66970 -6002
rect 52050 -6060 52110 -6026
rect 52430 -6059 52490 -6026
rect 52820 -6059 52880 -6026
rect 53200 -6059 53260 -6026
rect 52429 -6060 52490 -6059
rect 52620 -6060 52672 -6059
rect 52814 -6060 52880 -6059
rect 53198 -6060 53260 -6059
rect 53390 -6060 53442 -6059
rect 53580 -6060 53640 -6026
rect 53970 -6060 54030 -6026
rect 54350 -6060 54410 -6026
rect 54542 -6060 54594 -6059
rect 54740 -6060 54800 -6026
rect 55120 -6060 55180 -6026
rect 55310 -6060 55362 -6059
rect 55500 -6060 55560 -6026
rect 55890 -6059 55950 -6026
rect 55694 -6060 55746 -6059
rect 55886 -6060 55950 -6059
rect 56270 -6060 56330 -6026
rect 56462 -6060 56514 -6059
rect 56660 -6060 56720 -6026
rect 57040 -6060 57100 -6026
rect 57420 -6060 57480 -6026
rect 57810 -6059 57870 -6026
rect 57613 -6060 57665 -6059
rect 57804 -6060 57870 -6059
rect 58240 -6060 58300 -6026
rect 52050 -6061 57910 -6060
rect 49430 -6074 49482 -6064
rect 52047 -6069 57910 -6061
rect 52047 -6070 52429 -6069
rect 52047 -6071 52237 -6070
rect 49430 -6136 49482 -6126
rect 51842 -6120 51898 -6110
rect 49440 -6220 49470 -6136
rect 52099 -6092 52237 -6071
rect 52047 -6133 52099 -6123
rect 52289 -6092 52429 -6070
rect 52237 -6132 52289 -6122
rect 52481 -6092 52620 -6069
rect 52429 -6131 52481 -6121
rect 52672 -6092 52814 -6069
rect 52620 -6131 52672 -6121
rect 52866 -6070 53198 -6069
rect 52866 -6092 53004 -6070
rect 52814 -6131 52866 -6121
rect 53056 -6092 53198 -6070
rect 53004 -6132 53056 -6122
rect 53250 -6092 53390 -6069
rect 53198 -6131 53250 -6121
rect 53442 -6070 54542 -6069
rect 53442 -6092 53581 -6070
rect 53390 -6131 53442 -6121
rect 53633 -6092 53776 -6070
rect 53581 -6132 53633 -6122
rect 53828 -6092 53966 -6070
rect 53776 -6132 53828 -6122
rect 54018 -6092 54157 -6070
rect 53966 -6132 54018 -6122
rect 54209 -6092 54349 -6070
rect 54157 -6132 54209 -6122
rect 54401 -6092 54542 -6070
rect 54349 -6132 54401 -6122
rect 54594 -6070 55310 -6069
rect 54594 -6092 54734 -6070
rect 54542 -6131 54594 -6121
rect 54786 -6092 54926 -6070
rect 54734 -6132 54786 -6122
rect 54978 -6092 55119 -6070
rect 54926 -6132 54978 -6122
rect 55171 -6092 55310 -6070
rect 55119 -6132 55171 -6122
rect 55362 -6070 55694 -6069
rect 55362 -6092 55502 -6070
rect 55310 -6131 55362 -6121
rect 55554 -6092 55694 -6070
rect 55502 -6132 55554 -6122
rect 55746 -6092 55886 -6069
rect 55694 -6131 55746 -6121
rect 55938 -6070 56270 -6069
rect 55938 -6092 56077 -6070
rect 55886 -6131 55938 -6121
rect 56129 -6092 56270 -6070
rect 56077 -6132 56129 -6122
rect 56322 -6092 56462 -6069
rect 56270 -6131 56322 -6121
rect 56514 -6070 57613 -6069
rect 56514 -6092 56656 -6070
rect 56462 -6131 56514 -6121
rect 56708 -6071 57036 -6070
rect 56708 -6092 56847 -6071
rect 56656 -6132 56708 -6122
rect 56899 -6092 57036 -6071
rect 56847 -6133 56899 -6123
rect 57088 -6092 57229 -6070
rect 57036 -6132 57088 -6122
rect 57281 -6092 57422 -6070
rect 57229 -6132 57281 -6122
rect 57474 -6092 57613 -6070
rect 57422 -6132 57474 -6122
rect 57665 -6092 57804 -6069
rect 57613 -6131 57665 -6121
rect 57856 -6090 57910 -6069
rect 58100 -6061 58300 -6060
rect 58431 -6061 58483 -6059
rect 58620 -6061 58680 -6026
rect 59010 -6058 59070 -6026
rect 59400 -6058 59460 -6026
rect 58814 -6061 58866 -6058
rect 59008 -6061 59070 -6058
rect 59198 -6061 59250 -6059
rect 59392 -6061 59460 -6058
rect 59584 -6061 59636 -6058
rect 59780 -6059 59840 -6026
rect 59775 -6061 59840 -6059
rect 59970 -6061 60022 -6059
rect 60160 -6061 60220 -6026
rect 60351 -6061 60403 -6059
rect 60540 -6061 60600 -6026
rect 60736 -6061 60788 -6058
rect 60930 -6059 60990 -6026
rect 61320 -6059 61380 -6026
rect 60928 -6061 60990 -6059
rect 61120 -6061 61172 -6059
rect 61313 -6061 61380 -6059
rect 61504 -6061 61556 -6058
rect 61700 -6059 61760 -6026
rect 61696 -6061 61760 -6059
rect 61888 -6061 61940 -6058
rect 62080 -6061 62140 -6026
rect 62470 -6058 62530 -6026
rect 62271 -6061 62323 -6059
rect 62464 -6061 62530 -6058
rect 62656 -6061 62708 -6058
rect 62850 -6061 62910 -6026
rect 63041 -6061 63093 -6060
rect 63230 -6061 63290 -6026
rect 63620 -6059 63680 -6026
rect 64000 -6058 64060 -6026
rect 63423 -6061 63475 -6059
rect 63616 -6061 63680 -6059
rect 63807 -6061 63859 -6058
rect 63998 -6061 64060 -6058
rect 58100 -6068 64060 -6061
rect 58100 -6069 58623 -6068
rect 58100 -6070 58431 -6069
rect 58100 -6090 58241 -6070
rect 57804 -6131 57856 -6121
rect 58293 -6091 58431 -6070
rect 58241 -6132 58293 -6122
rect 58483 -6091 58623 -6069
rect 58431 -6131 58483 -6121
rect 58675 -6091 58814 -6068
rect 58623 -6130 58675 -6120
rect 58866 -6091 59008 -6068
rect 58814 -6130 58866 -6120
rect 59060 -6069 59392 -6068
rect 59060 -6091 59198 -6069
rect 59008 -6130 59060 -6120
rect 59250 -6091 59392 -6069
rect 59198 -6131 59250 -6121
rect 59444 -6091 59584 -6068
rect 59392 -6130 59444 -6120
rect 59636 -6069 60736 -6068
rect 59636 -6091 59775 -6069
rect 59584 -6130 59636 -6120
rect 59827 -6091 59970 -6069
rect 59775 -6131 59827 -6121
rect 60022 -6091 60160 -6069
rect 59970 -6131 60022 -6121
rect 60212 -6091 60351 -6069
rect 60160 -6131 60212 -6121
rect 60403 -6091 60543 -6069
rect 60351 -6131 60403 -6121
rect 60595 -6091 60736 -6069
rect 60543 -6131 60595 -6121
rect 60788 -6069 61504 -6068
rect 60788 -6091 60928 -6069
rect 60736 -6130 60788 -6120
rect 60980 -6091 61120 -6069
rect 60928 -6131 60980 -6121
rect 61172 -6091 61313 -6069
rect 61120 -6131 61172 -6121
rect 61365 -6091 61504 -6069
rect 61313 -6131 61365 -6121
rect 61556 -6069 61888 -6068
rect 61556 -6091 61696 -6069
rect 61504 -6130 61556 -6120
rect 61748 -6091 61888 -6069
rect 61696 -6131 61748 -6121
rect 61940 -6091 62080 -6068
rect 61888 -6130 61940 -6120
rect 62132 -6069 62464 -6068
rect 62132 -6091 62271 -6069
rect 62080 -6130 62132 -6120
rect 62323 -6091 62464 -6069
rect 62271 -6131 62323 -6121
rect 62516 -6091 62656 -6068
rect 62464 -6130 62516 -6120
rect 62708 -6069 63807 -6068
rect 62708 -6091 62850 -6069
rect 62656 -6130 62708 -6120
rect 62902 -6070 63230 -6069
rect 62902 -6091 63041 -6070
rect 62850 -6131 62902 -6121
rect 63093 -6091 63230 -6070
rect 63041 -6132 63093 -6122
rect 63282 -6091 63423 -6069
rect 63230 -6131 63282 -6121
rect 63475 -6091 63616 -6069
rect 63423 -6131 63475 -6121
rect 63668 -6091 63807 -6069
rect 63616 -6131 63668 -6121
rect 63859 -6091 63998 -6068
rect 63807 -6130 63859 -6120
rect 64050 -6070 64060 -6068
rect 63998 -6130 64050 -6120
rect 66930 -6142 66960 -6012
rect 51842 -6186 51898 -6176
rect 64128 -6176 64184 -6166
rect 49440 -6260 51556 -6220
rect 47224 -6678 47652 -6264
rect 51518 -6298 51556 -6260
rect 51516 -6308 51572 -6298
rect 51516 -6374 51572 -6364
rect 51726 -6382 51782 -6372
rect 51726 -6448 51782 -6438
rect 51726 -6552 51780 -6448
rect 51720 -6562 51780 -6552
rect 51776 -6612 51780 -6562
rect 51720 -6628 51776 -6618
rect 47224 -7752 47254 -6678
rect 47614 -7752 47652 -6678
rect 51842 -6680 51894 -6186
rect 51942 -6206 51998 -6196
rect 51942 -6272 51998 -6262
rect 52134 -6208 52190 -6198
rect 51942 -6288 51996 -6272
rect 52134 -6274 52190 -6264
rect 52328 -6210 52384 -6200
rect 51938 -6298 51996 -6288
rect 51994 -6334 51996 -6298
rect 51938 -6364 51994 -6354
rect 52136 -6424 52186 -6274
rect 52328 -6276 52384 -6266
rect 52524 -6210 52580 -6200
rect 52524 -6276 52580 -6266
rect 52714 -6214 52770 -6204
rect 52714 -6276 52770 -6270
rect 52906 -6210 52962 -6200
rect 52906 -6276 52962 -6266
rect 53100 -6212 53156 -6202
rect 52330 -6288 52384 -6276
rect 52330 -6298 52386 -6288
rect 52330 -6364 52386 -6354
rect 52528 -6422 52578 -6276
rect 52714 -6280 52772 -6276
rect 52716 -6286 52772 -6280
rect 52716 -6352 52772 -6342
rect 52910 -6422 52960 -6276
rect 53100 -6278 53156 -6268
rect 53288 -6210 53344 -6200
rect 53288 -6270 53344 -6266
rect 53480 -6212 53536 -6202
rect 53672 -6208 53728 -6198
rect 53536 -6268 53540 -6230
rect 53288 -6276 53350 -6270
rect 53102 -6288 53158 -6278
rect 53102 -6354 53158 -6344
rect 52132 -6434 52188 -6424
rect 52132 -6500 52188 -6490
rect 52510 -6432 52578 -6422
rect 52566 -6456 52578 -6432
rect 52908 -6432 52964 -6422
rect 53300 -6424 53350 -6276
rect 53480 -6278 53540 -6268
rect 53672 -6274 53728 -6264
rect 53870 -6210 53926 -6200
rect 53486 -6286 53540 -6278
rect 53486 -6296 53542 -6286
rect 53486 -6362 53542 -6352
rect 53676 -6424 53726 -6274
rect 53870 -6276 53926 -6266
rect 53872 -6284 53926 -6276
rect 54058 -6212 54114 -6202
rect 54058 -6278 54114 -6268
rect 54252 -6210 54308 -6200
rect 54440 -6208 54496 -6198
rect 54308 -6266 54310 -6230
rect 54252 -6276 54310 -6266
rect 53872 -6294 53928 -6284
rect 53872 -6360 53928 -6350
rect 52510 -6498 52566 -6488
rect 52908 -6498 52964 -6488
rect 53294 -6434 53350 -6424
rect 53294 -6500 53350 -6490
rect 53672 -6434 53728 -6424
rect 54064 -6426 54114 -6278
rect 54256 -6286 54310 -6276
rect 54438 -6264 54440 -6262
rect 54438 -6274 54496 -6264
rect 54632 -6214 54688 -6204
rect 54826 -6212 54882 -6202
rect 54688 -6270 54692 -6238
rect 54256 -6296 54312 -6286
rect 54256 -6362 54312 -6352
rect 54438 -6426 54488 -6274
rect 54632 -6280 54692 -6270
rect 54638 -6288 54692 -6280
rect 54824 -6268 54826 -6264
rect 54824 -6278 54882 -6268
rect 55016 -6212 55072 -6202
rect 55212 -6212 55268 -6202
rect 55016 -6278 55072 -6268
rect 54638 -6298 54694 -6288
rect 54638 -6364 54694 -6354
rect 54824 -6426 54874 -6278
rect 55018 -6282 55072 -6278
rect 55202 -6268 55212 -6262
rect 55202 -6278 55268 -6268
rect 55402 -6212 55458 -6202
rect 55594 -6210 55650 -6200
rect 55458 -6268 55466 -6232
rect 55402 -6278 55466 -6268
rect 55786 -6208 55842 -6198
rect 55594 -6276 55650 -6266
rect 55784 -6264 55786 -6232
rect 55784 -6274 55842 -6264
rect 55978 -6210 56034 -6200
rect 55018 -6292 55074 -6282
rect 55018 -6358 55074 -6348
rect 55202 -6426 55252 -6278
rect 55412 -6294 55466 -6278
rect 55412 -6304 55468 -6294
rect 55412 -6370 55468 -6360
rect 55598 -6422 55648 -6276
rect 55784 -6292 55838 -6274
rect 55782 -6302 55838 -6292
rect 55782 -6368 55838 -6358
rect 55978 -6276 56034 -6266
rect 56172 -6208 56228 -6198
rect 56362 -6212 56418 -6202
rect 56172 -6274 56228 -6264
rect 53672 -6500 53728 -6490
rect 54056 -6436 54114 -6426
rect 54112 -6460 54114 -6436
rect 54428 -6436 54488 -6426
rect 54056 -6502 54112 -6492
rect 54484 -6450 54488 -6436
rect 54820 -6436 54876 -6426
rect 54428 -6502 54484 -6492
rect 54820 -6502 54876 -6492
rect 55198 -6436 55254 -6426
rect 55198 -6502 55254 -6492
rect 55594 -6432 55650 -6422
rect 55978 -6424 56028 -6276
rect 56174 -6288 56228 -6274
rect 56360 -6268 56362 -6260
rect 56360 -6278 56418 -6268
rect 56558 -6210 56614 -6200
rect 56558 -6276 56614 -6266
rect 56746 -6210 56802 -6200
rect 56940 -6210 56996 -6200
rect 56746 -6276 56802 -6266
rect 56174 -6298 56230 -6288
rect 56174 -6364 56230 -6354
rect 55594 -6498 55650 -6488
rect 55974 -6434 56030 -6424
rect 56360 -6426 56410 -6278
rect 56560 -6290 56614 -6276
rect 56560 -6300 56616 -6290
rect 56560 -6366 56616 -6356
rect 56752 -6426 56802 -6276
rect 56938 -6266 56940 -6232
rect 57132 -6210 57188 -6200
rect 56938 -6276 56996 -6266
rect 57130 -6266 57132 -6256
rect 57318 -6214 57374 -6204
rect 57130 -6276 57188 -6266
rect 57314 -6270 57318 -6240
rect 57516 -6212 57572 -6202
rect 56938 -6286 56992 -6276
rect 56936 -6296 56992 -6286
rect 56936 -6362 56992 -6352
rect 57130 -6426 57180 -6276
rect 57314 -6280 57374 -6270
rect 57506 -6268 57516 -6254
rect 57506 -6278 57572 -6268
rect 57702 -6212 57758 -6202
rect 58138 -6210 58194 -6200
rect 57758 -6268 57762 -6240
rect 57702 -6278 57762 -6268
rect 57314 -6290 57368 -6280
rect 57312 -6300 57368 -6290
rect 57312 -6366 57368 -6356
rect 57506 -6426 57556 -6278
rect 57708 -6288 57762 -6278
rect 58130 -6266 58138 -6238
rect 58330 -6212 58386 -6202
rect 58130 -6276 58194 -6266
rect 58326 -6268 58330 -6254
rect 58526 -6210 58582 -6200
rect 58130 -6282 58184 -6276
rect 57708 -6298 57764 -6288
rect 57708 -6364 57764 -6354
rect 58128 -6292 58184 -6282
rect 58128 -6358 58184 -6348
rect 58326 -6278 58386 -6268
rect 58522 -6266 58526 -6240
rect 58522 -6276 58582 -6266
rect 58714 -6212 58770 -6202
rect 58326 -6426 58376 -6278
rect 58522 -6284 58576 -6276
rect 58714 -6278 58770 -6268
rect 58906 -6214 58962 -6204
rect 58520 -6294 58576 -6284
rect 58520 -6360 58576 -6350
rect 58716 -6426 58766 -6278
rect 58906 -6280 58962 -6270
rect 58908 -6284 58962 -6280
rect 59100 -6212 59156 -6202
rect 59100 -6278 59156 -6268
rect 59292 -6214 59348 -6204
rect 58908 -6294 58964 -6284
rect 58908 -6360 58964 -6350
rect 59100 -6424 59150 -6278
rect 59292 -6280 59348 -6270
rect 59484 -6212 59540 -6202
rect 59678 -6210 59734 -6200
rect 59540 -6268 59542 -6258
rect 59484 -6278 59542 -6268
rect 59868 -6210 59924 -6200
rect 59734 -6266 59744 -6242
rect 59678 -6276 59744 -6266
rect 59292 -6288 59346 -6280
rect 59290 -6298 59346 -6288
rect 59290 -6364 59346 -6354
rect 55974 -6500 56030 -6490
rect 56352 -6436 56410 -6426
rect 56408 -6448 56410 -6436
rect 56744 -6436 56802 -6426
rect 56352 -6502 56408 -6492
rect 56800 -6448 56802 -6436
rect 57126 -6436 57182 -6426
rect 56744 -6502 56800 -6492
rect 57126 -6502 57182 -6492
rect 57500 -6436 57556 -6426
rect 57500 -6502 57556 -6492
rect 58322 -6436 58378 -6426
rect 58322 -6502 58378 -6492
rect 58712 -6436 58768 -6426
rect 58712 -6502 58768 -6492
rect 59100 -6434 59156 -6424
rect 59492 -6426 59542 -6278
rect 59690 -6286 59744 -6276
rect 59862 -6266 59868 -6256
rect 59862 -6276 59924 -6266
rect 60060 -6214 60116 -6204
rect 60252 -6214 60308 -6204
rect 60116 -6270 60120 -6232
rect 59690 -6296 59746 -6286
rect 59690 -6362 59746 -6352
rect 59862 -6426 59912 -6276
rect 60060 -6280 60120 -6270
rect 60444 -6212 60500 -6202
rect 60252 -6280 60308 -6270
rect 60440 -6268 60444 -6244
rect 60440 -6278 60500 -6268
rect 60638 -6212 60694 -6202
rect 60828 -6214 60884 -6204
rect 60694 -6268 60696 -6258
rect 60638 -6278 60696 -6268
rect 60066 -6290 60122 -6280
rect 60066 -6356 60122 -6346
rect 60256 -6426 60306 -6280
rect 60440 -6284 60494 -6278
rect 60438 -6294 60494 -6284
rect 60438 -6360 60494 -6350
rect 60646 -6424 60696 -6278
rect 61018 -6212 61074 -6202
rect 60884 -6270 60890 -6240
rect 60828 -6280 60890 -6270
rect 60836 -6290 60890 -6280
rect 61018 -6278 61074 -6268
rect 61212 -6208 61268 -6198
rect 61404 -6214 61460 -6204
rect 61268 -6264 61272 -6244
rect 61212 -6274 61272 -6264
rect 60836 -6300 60892 -6290
rect 60836 -6366 60892 -6356
rect 61018 -6424 61068 -6278
rect 61218 -6286 61272 -6274
rect 61596 -6214 61652 -6204
rect 61404 -6280 61460 -6270
rect 61218 -6296 61274 -6286
rect 61218 -6362 61274 -6352
rect 61410 -6422 61460 -6280
rect 61594 -6270 61596 -6234
rect 61594 -6280 61652 -6270
rect 61786 -6214 61842 -6204
rect 61976 -6212 62032 -6202
rect 61786 -6280 61842 -6270
rect 61974 -6268 61976 -6238
rect 62174 -6210 62230 -6200
rect 61974 -6278 62032 -6268
rect 62170 -6266 62174 -6262
rect 62364 -6214 62420 -6204
rect 62170 -6276 62230 -6266
rect 62362 -6270 62364 -6236
rect 61594 -6284 61648 -6280
rect 61592 -6294 61648 -6284
rect 61592 -6360 61648 -6350
rect 59100 -6500 59156 -6490
rect 59490 -6436 59546 -6426
rect 59490 -6502 59546 -6492
rect 59858 -6436 59914 -6426
rect 59858 -6502 59914 -6492
rect 60252 -6436 60308 -6426
rect 60252 -6502 60308 -6492
rect 60644 -6434 60700 -6424
rect 60644 -6500 60700 -6490
rect 61010 -6434 61068 -6424
rect 61066 -6446 61068 -6434
rect 61406 -6432 61462 -6422
rect 61786 -6426 61836 -6280
rect 61974 -6286 62028 -6278
rect 61972 -6296 62028 -6286
rect 61972 -6362 62028 -6352
rect 62170 -6424 62220 -6276
rect 62362 -6280 62420 -6270
rect 62554 -6212 62610 -6202
rect 62750 -6212 62806 -6202
rect 62554 -6278 62610 -6268
rect 62744 -6268 62750 -6242
rect 62744 -6278 62806 -6268
rect 62938 -6210 62994 -6200
rect 63134 -6214 63190 -6204
rect 62938 -6276 62994 -6266
rect 63130 -6270 63134 -6238
rect 63322 -6212 63378 -6202
rect 62362 -6286 62416 -6280
rect 62360 -6296 62416 -6286
rect 62360 -6362 62416 -6352
rect 61010 -6500 61066 -6490
rect 61406 -6498 61462 -6488
rect 61782 -6436 61838 -6426
rect 61782 -6502 61838 -6492
rect 62162 -6434 62220 -6424
rect 62556 -6426 62606 -6278
rect 62744 -6284 62798 -6278
rect 62742 -6294 62798 -6284
rect 62742 -6360 62798 -6350
rect 62942 -6424 62992 -6276
rect 63130 -6280 63190 -6270
rect 63320 -6268 63322 -6256
rect 63320 -6278 63378 -6268
rect 63512 -6210 63568 -6200
rect 63512 -6276 63568 -6266
rect 63710 -6212 63766 -6202
rect 63902 -6210 63958 -6200
rect 63130 -6286 63184 -6280
rect 63128 -6296 63184 -6286
rect 63128 -6362 63184 -6352
rect 62218 -6450 62220 -6434
rect 62550 -6436 62606 -6426
rect 62162 -6500 62218 -6490
rect 62550 -6502 62606 -6492
rect 62936 -6434 62992 -6424
rect 63320 -6426 63370 -6278
rect 63512 -6284 63566 -6276
rect 63510 -6294 63566 -6284
rect 63510 -6360 63566 -6350
rect 63710 -6278 63766 -6268
rect 63900 -6266 63902 -6242
rect 64528 -6172 66960 -6142
rect 64184 -6232 64196 -6216
rect 64128 -6242 64196 -6232
rect 63900 -6276 63958 -6266
rect 63710 -6424 63760 -6278
rect 63900 -6282 63954 -6276
rect 63898 -6292 63954 -6282
rect 63898 -6358 63954 -6348
rect 62936 -6500 62992 -6490
rect 63316 -6436 63372 -6426
rect 63316 -6502 63372 -6492
rect 63706 -6434 63762 -6424
rect 63706 -6500 63762 -6490
rect 52238 -6562 52294 -6552
rect 52236 -6618 52238 -6606
rect 52620 -6562 52676 -6552
rect 52294 -6618 52298 -6606
rect 49440 -6690 51894 -6680
rect 49440 -6720 51838 -6690
rect 49440 -6862 49470 -6720
rect 51838 -6756 51894 -6746
rect 52044 -6690 52100 -6680
rect 52236 -6690 52298 -6618
rect 52618 -6618 52620 -6604
rect 53002 -6562 53058 -6552
rect 52676 -6618 52680 -6604
rect 52236 -6724 52238 -6690
rect 52044 -6756 52100 -6746
rect 52294 -6724 52298 -6690
rect 52432 -6696 52488 -6686
rect 52238 -6756 52294 -6746
rect 52618 -6692 52680 -6618
rect 53390 -6562 53446 -6552
rect 53058 -6618 53064 -6608
rect 52618 -6722 52622 -6692
rect 52432 -6762 52488 -6752
rect 52678 -6722 52680 -6692
rect 52818 -6692 52874 -6682
rect 52622 -6758 52678 -6748
rect 53002 -6692 53064 -6618
rect 53768 -6562 53824 -6552
rect 53446 -6618 53452 -6604
rect 53002 -6726 53006 -6692
rect 52818 -6758 52874 -6748
rect 53062 -6726 53064 -6692
rect 53200 -6690 53256 -6680
rect 53006 -6758 53062 -6748
rect 53390 -6690 53452 -6618
rect 54150 -6562 54206 -6552
rect 53824 -6618 53830 -6604
rect 53390 -6722 53394 -6690
rect 53200 -6756 53256 -6746
rect 53450 -6722 53452 -6690
rect 53582 -6692 53638 -6682
rect 53394 -6756 53450 -6746
rect 53768 -6690 53830 -6618
rect 54538 -6562 54594 -6552
rect 54206 -6618 54212 -6604
rect 53768 -6722 53774 -6690
rect 53582 -6758 53638 -6748
rect 53774 -6756 53830 -6746
rect 53964 -6694 54020 -6684
rect 54150 -6692 54212 -6618
rect 54920 -6562 54976 -6552
rect 54594 -6618 54600 -6602
rect 54150 -6722 54156 -6692
rect 53964 -6760 54020 -6750
rect 54156 -6758 54212 -6748
rect 54350 -6694 54406 -6684
rect 54538 -6690 54600 -6618
rect 55304 -6562 55360 -6552
rect 54976 -6618 54982 -6604
rect 54538 -6720 54542 -6690
rect 54350 -6760 54406 -6750
rect 54598 -6720 54600 -6690
rect 54740 -6692 54796 -6682
rect 54542 -6756 54598 -6746
rect 54920 -6690 54982 -6618
rect 55682 -6562 55738 -6552
rect 55360 -6618 55366 -6602
rect 54920 -6722 54926 -6690
rect 54740 -6758 54796 -6748
rect 54926 -6756 54982 -6746
rect 55120 -6696 55176 -6686
rect 55304 -6692 55366 -6618
rect 56072 -6562 56128 -6552
rect 55738 -6618 55744 -6602
rect 55682 -6680 55744 -6618
rect 56454 -6562 56510 -6552
rect 56128 -6618 56134 -6598
rect 55304 -6720 55310 -6692
rect 55120 -6762 55176 -6752
rect 55310 -6758 55366 -6748
rect 55502 -6696 55558 -6686
rect 55682 -6690 55746 -6680
rect 55682 -6720 55690 -6690
rect 55502 -6762 55558 -6752
rect 55690 -6756 55746 -6746
rect 55886 -6694 55942 -6684
rect 56072 -6688 56134 -6618
rect 56840 -6562 56896 -6552
rect 56510 -6618 56516 -6606
rect 56072 -6716 56078 -6688
rect 55886 -6760 55942 -6750
rect 56078 -6754 56134 -6744
rect 56272 -6692 56328 -6682
rect 56454 -6694 56516 -6618
rect 57222 -6562 57278 -6552
rect 56896 -6618 56902 -6600
rect 56840 -6680 56902 -6618
rect 57602 -6562 57658 -6552
rect 57278 -6618 57284 -6602
rect 56454 -6724 56460 -6694
rect 56272 -6758 56328 -6748
rect 56460 -6760 56516 -6750
rect 56658 -6694 56714 -6684
rect 56840 -6690 56904 -6680
rect 56840 -6718 56848 -6690
rect 56658 -6760 56714 -6750
rect 56848 -6756 56904 -6746
rect 57038 -6696 57094 -6686
rect 57222 -6690 57284 -6618
rect 58414 -6562 58470 -6552
rect 57658 -6618 57664 -6602
rect 57222 -6720 57228 -6690
rect 57038 -6762 57094 -6752
rect 57228 -6756 57284 -6746
rect 57422 -6696 57478 -6686
rect 57602 -6692 57664 -6618
rect 58412 -6618 58414 -6600
rect 58796 -6562 58852 -6552
rect 58470 -6618 58474 -6600
rect 58412 -6682 58474 -6618
rect 59186 -6562 59242 -6552
rect 58852 -6618 58858 -6600
rect 57602 -6720 57608 -6692
rect 57422 -6762 57478 -6752
rect 57608 -6758 57664 -6748
rect 57806 -6694 57862 -6684
rect 57806 -6760 57862 -6750
rect 58230 -6694 58286 -6684
rect 58412 -6692 58476 -6682
rect 58412 -6718 58420 -6692
rect 58230 -6760 58286 -6750
rect 58420 -6758 58476 -6748
rect 58612 -6698 58668 -6688
rect 58796 -6692 58858 -6618
rect 59568 -6562 59624 -6552
rect 59242 -6618 59248 -6600
rect 58796 -6718 58802 -6692
rect 58612 -6764 58668 -6754
rect 58802 -6758 58858 -6748
rect 58996 -6694 59052 -6684
rect 59186 -6690 59248 -6618
rect 59566 -6618 59568 -6600
rect 59954 -6562 60010 -6552
rect 59624 -6618 59628 -6600
rect 59186 -6718 59190 -6690
rect 58996 -6760 59052 -6750
rect 59246 -6718 59248 -6690
rect 59382 -6694 59438 -6684
rect 59190 -6756 59246 -6746
rect 59566 -6692 59628 -6618
rect 60336 -6562 60392 -6552
rect 60010 -6618 60018 -6598
rect 59954 -6628 60018 -6618
rect 59566 -6718 59572 -6692
rect 59382 -6760 59438 -6750
rect 59572 -6758 59628 -6748
rect 59764 -6694 59820 -6684
rect 59956 -6690 60018 -6628
rect 60722 -6562 60778 -6552
rect 60392 -6618 60398 -6600
rect 59956 -6716 59960 -6690
rect 59764 -6760 59820 -6750
rect 60016 -6716 60018 -6690
rect 60154 -6692 60210 -6682
rect 59960 -6756 60016 -6746
rect 60336 -6690 60398 -6618
rect 61104 -6562 61160 -6552
rect 60778 -6618 60784 -6600
rect 60336 -6718 60342 -6690
rect 60154 -6758 60210 -6748
rect 60342 -6756 60398 -6746
rect 60534 -6696 60590 -6686
rect 60722 -6688 60784 -6618
rect 61482 -6562 61538 -6552
rect 61160 -6618 61166 -6602
rect 60722 -6718 60726 -6688
rect 60534 -6762 60590 -6752
rect 60782 -6718 60784 -6688
rect 60918 -6694 60974 -6684
rect 60726 -6754 60782 -6744
rect 61104 -6690 61166 -6618
rect 61866 -6562 61922 -6552
rect 61538 -6618 61546 -6602
rect 61482 -6628 61546 -6618
rect 61484 -6680 61546 -6628
rect 62252 -6562 62308 -6552
rect 61922 -6618 61928 -6602
rect 61866 -6680 61928 -6618
rect 62640 -6562 62696 -6552
rect 62308 -6618 62314 -6602
rect 62252 -6680 62314 -6618
rect 62638 -6618 62640 -6600
rect 63022 -6562 63078 -6552
rect 62696 -6618 62700 -6600
rect 61104 -6720 61110 -6690
rect 60918 -6760 60974 -6750
rect 61110 -6756 61166 -6746
rect 61300 -6694 61356 -6684
rect 61484 -6690 61548 -6680
rect 61484 -6720 61492 -6690
rect 61300 -6760 61356 -6750
rect 61492 -6756 61548 -6746
rect 61688 -6696 61744 -6686
rect 61866 -6690 61930 -6680
rect 61866 -6720 61874 -6690
rect 61688 -6762 61744 -6752
rect 61874 -6756 61930 -6746
rect 62070 -6692 62126 -6682
rect 62252 -6690 62316 -6680
rect 62252 -6720 62260 -6690
rect 62070 -6758 62126 -6748
rect 62260 -6756 62316 -6746
rect 62456 -6692 62512 -6682
rect 62638 -6690 62700 -6618
rect 63406 -6562 63462 -6552
rect 63078 -6618 63084 -6602
rect 62638 -6718 62644 -6690
rect 62456 -6758 62512 -6748
rect 62644 -6756 62700 -6746
rect 62840 -6690 62896 -6680
rect 63022 -6692 63084 -6618
rect 63792 -6562 63848 -6552
rect 63462 -6618 63468 -6602
rect 63022 -6720 63028 -6692
rect 62840 -6756 62896 -6746
rect 63028 -6758 63084 -6748
rect 63220 -6692 63276 -6682
rect 63406 -6692 63468 -6618
rect 63848 -6618 63854 -6600
rect 63406 -6720 63412 -6692
rect 63220 -6758 63276 -6748
rect 63412 -6758 63468 -6748
rect 63608 -6690 63664 -6680
rect 63792 -6688 63854 -6618
rect 64144 -6680 64196 -6242
rect 64236 -6400 64292 -6390
rect 64528 -6426 64562 -6172
rect 64236 -6466 64292 -6456
rect 64502 -6436 64562 -6426
rect 64236 -6552 64288 -6466
rect 64558 -6484 64562 -6436
rect 68894 -6272 68930 -5188
rect 69296 -6272 69326 -5188
rect 64502 -6502 64558 -6492
rect 64236 -6562 64294 -6552
rect 64236 -6608 64238 -6562
rect 64294 -6618 64558 -6582
rect 64238 -6620 64558 -6618
rect 64238 -6628 64294 -6620
rect 64530 -6680 64558 -6620
rect 68894 -6672 69326 -6272
rect 63792 -6718 63796 -6688
rect 63608 -6756 63664 -6746
rect 63852 -6718 63854 -6688
rect 63992 -6690 64048 -6680
rect 63796 -6754 63852 -6744
rect 63992 -6756 64048 -6746
rect 64144 -6690 64200 -6680
rect 64530 -6710 66950 -6680
rect 64144 -6756 64200 -6746
rect 51950 -6826 63950 -6810
rect 51950 -6827 59100 -6826
rect 51950 -6828 52912 -6827
rect 49436 -6872 49488 -6862
rect 52002 -6880 52142 -6828
rect 52194 -6880 52335 -6828
rect 52387 -6880 52527 -6828
rect 52579 -6880 52720 -6828
rect 52772 -6879 52912 -6828
rect 52964 -6828 53487 -6827
rect 52964 -6879 53103 -6828
rect 52772 -6880 53103 -6879
rect 53155 -6880 53295 -6828
rect 53347 -6879 53487 -6828
rect 53539 -6879 53679 -6827
rect 53731 -6828 54063 -6827
rect 53731 -6879 53871 -6828
rect 53347 -6880 53871 -6879
rect 53923 -6879 54063 -6828
rect 54115 -6828 54446 -6827
rect 54115 -6879 54255 -6828
rect 53923 -6880 54255 -6879
rect 54307 -6879 54446 -6828
rect 54498 -6828 55599 -6827
rect 54498 -6879 54640 -6828
rect 54307 -6880 54640 -6879
rect 54692 -6880 54830 -6828
rect 54882 -6880 55022 -6828
rect 55074 -6880 55215 -6828
rect 55267 -6880 55406 -6828
rect 55458 -6879 55599 -6828
rect 55651 -6828 56560 -6827
rect 55651 -6879 55792 -6828
rect 55458 -6880 55792 -6879
rect 55844 -6880 55983 -6828
rect 56035 -6880 56176 -6828
rect 56228 -6880 56366 -6828
rect 56418 -6879 56560 -6828
rect 56612 -6828 57518 -6827
rect 56612 -6879 56749 -6828
rect 56418 -6880 56749 -6879
rect 56801 -6880 56942 -6828
rect 56994 -6880 57135 -6828
rect 57187 -6880 57325 -6828
rect 57377 -6879 57518 -6828
rect 57570 -6879 57707 -6827
rect 57759 -6879 58138 -6827
rect 58190 -6879 58330 -6827
rect 58382 -6879 58523 -6827
rect 58575 -6879 58715 -6827
rect 58767 -6879 58908 -6827
rect 58960 -6878 59100 -6827
rect 59152 -6827 59675 -6826
rect 59152 -6878 59291 -6827
rect 58960 -6879 59291 -6878
rect 59343 -6879 59483 -6827
rect 59535 -6878 59675 -6827
rect 59727 -6878 59867 -6826
rect 59919 -6827 60251 -6826
rect 59919 -6878 60059 -6827
rect 59535 -6879 60059 -6878
rect 60111 -6878 60251 -6827
rect 60303 -6827 60634 -6826
rect 60303 -6878 60443 -6827
rect 60111 -6879 60443 -6878
rect 60495 -6878 60634 -6827
rect 60686 -6827 61787 -6826
rect 60686 -6878 60828 -6827
rect 60495 -6879 60828 -6878
rect 60880 -6879 61018 -6827
rect 61070 -6879 61210 -6827
rect 61262 -6879 61403 -6827
rect 61455 -6879 61594 -6827
rect 61646 -6878 61787 -6827
rect 61839 -6827 62748 -6826
rect 61839 -6878 61980 -6827
rect 61646 -6879 61980 -6878
rect 62032 -6879 62171 -6827
rect 62223 -6879 62364 -6827
rect 62416 -6879 62554 -6827
rect 62606 -6878 62748 -6827
rect 62800 -6827 63706 -6826
rect 62800 -6878 62937 -6827
rect 62606 -6879 62937 -6878
rect 62989 -6879 63130 -6827
rect 63182 -6879 63323 -6827
rect 63375 -6879 63513 -6827
rect 63565 -6878 63706 -6827
rect 63758 -6878 63895 -6826
rect 63947 -6878 63950 -6826
rect 66920 -6840 66950 -6710
rect 63565 -6879 63950 -6878
rect 57377 -6880 63950 -6879
rect 51950 -6890 63950 -6880
rect 66912 -6850 66964 -6840
rect 49436 -6934 49488 -6924
rect 52000 -7040 52060 -6890
rect 52390 -7040 52450 -6890
rect 52960 -7040 53020 -6890
rect 53350 -7040 53410 -6890
rect 53730 -7040 53790 -6890
rect 54120 -7040 54180 -6890
rect 54510 -7040 54570 -6890
rect 54890 -7040 54950 -6890
rect 55260 -7040 55320 -6890
rect 55650 -7040 55710 -6890
rect 56030 -7040 56090 -6890
rect 56410 -7040 56470 -6890
rect 56810 -7040 56870 -6890
rect 57180 -7040 57240 -6890
rect 57570 -7040 57630 -6890
rect 57960 -7040 58020 -6890
rect 58340 -7040 58400 -6890
rect 58730 -7040 58790 -6890
rect 59110 -7040 59170 -6890
rect 59490 -7040 59550 -6890
rect 59880 -7040 59940 -6890
rect 60260 -7040 60320 -6890
rect 60640 -7040 60700 -6890
rect 61030 -7040 61090 -6890
rect 61420 -7040 61480 -6890
rect 61800 -7040 61860 -6890
rect 62180 -7040 62240 -6890
rect 62570 -7040 62630 -6890
rect 62950 -7040 63010 -6890
rect 63340 -7040 63400 -6890
rect 63720 -7040 63780 -6890
rect 66912 -6912 66964 -6902
rect 51992 -7112 63790 -7040
rect 50087 -7300 50139 -7292
rect 50277 -7300 50329 -7291
rect 50470 -7300 50522 -7294
rect 50662 -7299 50714 -7289
rect 50087 -7301 50662 -7300
rect 50087 -7302 50277 -7301
rect 50139 -7330 50277 -7302
rect 50087 -7364 50139 -7354
rect 50329 -7304 50662 -7301
rect 50329 -7330 50470 -7304
rect 50277 -7363 50329 -7353
rect 50522 -7330 50662 -7304
rect 50470 -7366 50522 -7356
rect 50854 -7300 50906 -7293
rect 51046 -7298 51098 -7288
rect 50714 -7303 51046 -7300
rect 50714 -7330 50854 -7303
rect 50662 -7361 50714 -7351
rect 50906 -7330 51046 -7303
rect 50854 -7365 50906 -7355
rect 51238 -7299 51290 -7289
rect 51098 -7330 51238 -7300
rect 51046 -7360 51098 -7350
rect 51428 -7298 51480 -7288
rect 51290 -7330 51428 -7300
rect 51238 -7361 51290 -7351
rect 51622 -7300 51674 -7299
rect 51811 -7300 51863 -7297
rect 52000 -7300 52060 -7112
rect 52200 -7300 52252 -7298
rect 52390 -7300 52450 -7112
rect 52582 -7300 52634 -7298
rect 52774 -7300 52826 -7291
rect 52960 -7300 53020 -7112
rect 53159 -7300 53211 -7292
rect 53350 -7300 53410 -7112
rect 53542 -7300 53594 -7290
rect 53730 -7300 53790 -7112
rect 54120 -7287 54180 -7112
rect 53927 -7300 53979 -7291
rect 54119 -7297 54180 -7287
rect 54510 -7291 54570 -7112
rect 54890 -7290 54950 -7112
rect 55260 -7288 55320 -7112
rect 51480 -7301 53351 -7300
rect 51480 -7307 52774 -7301
rect 51480 -7309 51811 -7307
rect 51480 -7330 51622 -7309
rect 51428 -7360 51480 -7350
rect 51674 -7330 51811 -7309
rect 51622 -7371 51674 -7361
rect 51863 -7330 52001 -7307
rect 51811 -7369 51863 -7359
rect 52053 -7308 52392 -7307
rect 52053 -7330 52200 -7308
rect 52001 -7369 52053 -7359
rect 52252 -7330 52392 -7308
rect 52200 -7370 52252 -7360
rect 52444 -7308 52774 -7307
rect 52444 -7330 52582 -7308
rect 52392 -7369 52444 -7359
rect 52634 -7330 52774 -7308
rect 52582 -7370 52634 -7360
rect 52826 -7302 53351 -7301
rect 52826 -7303 53159 -7302
rect 52826 -7330 52966 -7303
rect 52774 -7363 52826 -7353
rect 53018 -7330 53159 -7303
rect 52966 -7365 53018 -7355
rect 53211 -7330 53351 -7302
rect 53159 -7364 53211 -7354
rect 53403 -7330 53542 -7300
rect 53351 -7362 53403 -7352
rect 53594 -7301 54119 -7300
rect 53594 -7305 53927 -7301
rect 53594 -7330 53736 -7305
rect 53542 -7362 53594 -7352
rect 53788 -7330 53927 -7305
rect 53736 -7367 53788 -7357
rect 53979 -7330 54119 -7301
rect 53927 -7363 53979 -7353
rect 54171 -7300 54180 -7297
rect 54312 -7300 54364 -7291
rect 54504 -7300 54570 -7291
rect 54697 -7300 54749 -7292
rect 54889 -7300 54950 -7290
rect 55080 -7299 55132 -7289
rect 54171 -7301 54889 -7300
rect 54171 -7330 54312 -7301
rect 54119 -7359 54171 -7349
rect 54364 -7330 54504 -7301
rect 54312 -7363 54364 -7353
rect 54556 -7302 54889 -7301
rect 54556 -7330 54697 -7302
rect 54504 -7363 54556 -7353
rect 54749 -7330 54889 -7302
rect 54697 -7364 54749 -7354
rect 54941 -7330 55080 -7300
rect 54889 -7362 54941 -7352
rect 55260 -7298 55323 -7288
rect 55260 -7300 55271 -7298
rect 55132 -7330 55271 -7300
rect 55080 -7361 55132 -7351
rect 55464 -7298 55516 -7288
rect 55323 -7330 55464 -7300
rect 55271 -7360 55323 -7350
rect 55650 -7300 55710 -7112
rect 55846 -7300 55898 -7298
rect 56030 -7300 56090 -7112
rect 56410 -7300 56470 -7112
rect 56810 -7300 56870 -7112
rect 57180 -7296 57240 -7112
rect 56997 -7300 57049 -7298
rect 57180 -7300 57243 -7296
rect 57384 -7300 57436 -7297
rect 57570 -7300 57630 -7112
rect 57960 -7298 58020 -7112
rect 57766 -7300 57818 -7298
rect 57959 -7300 58020 -7298
rect 58151 -7300 58203 -7298
rect 58340 -7300 58400 -7112
rect 58730 -7297 58790 -7112
rect 58535 -7300 58587 -7298
rect 58726 -7300 58790 -7297
rect 58921 -7300 58973 -7298
rect 59110 -7300 59170 -7112
rect 59303 -7300 59355 -7298
rect 59490 -7300 59550 -7112
rect 59880 -7298 59940 -7112
rect 59686 -7300 59738 -7298
rect 59878 -7300 59940 -7298
rect 60071 -7300 60123 -7298
rect 60260 -7300 60320 -7112
rect 60454 -7300 60506 -7298
rect 60640 -7300 60700 -7112
rect 60838 -7300 60890 -7298
rect 61030 -7300 61090 -7112
rect 61420 -7297 61480 -7112
rect 61222 -7300 61274 -7299
rect 61415 -7300 61480 -7297
rect 61605 -7300 61657 -7297
rect 61800 -7299 61860 -7112
rect 61798 -7300 61860 -7299
rect 61990 -7300 62042 -7298
rect 62180 -7300 62240 -7112
rect 62374 -7300 62426 -7297
rect 62570 -7298 62630 -7112
rect 62950 -7298 63010 -7112
rect 62566 -7300 62630 -7298
rect 62757 -7300 62809 -7298
rect 62949 -7300 63010 -7298
rect 63143 -7300 63195 -7297
rect 63340 -7298 63400 -7112
rect 63335 -7300 63400 -7298
rect 63525 -7300 63577 -7299
rect 63720 -7300 63780 -7112
rect 63909 -7300 63961 -7298
rect 64102 -7300 64154 -7297
rect 64295 -7300 64347 -7298
rect 64486 -7300 64538 -7298
rect 64677 -7300 64729 -7298
rect 64870 -7300 64922 -7298
rect 65063 -7300 65115 -7298
rect 65254 -7300 65306 -7298
rect 65445 -7300 65497 -7297
rect 65636 -7300 65688 -7297
rect 65829 -7300 65881 -7298
rect 66023 -7300 66075 -7298
rect 66211 -7300 66263 -7299
rect 55516 -7306 66470 -7300
rect 55516 -7307 57191 -7306
rect 55516 -7330 55655 -7307
rect 55464 -7360 55516 -7350
rect 55707 -7308 57191 -7307
rect 55707 -7330 55846 -7308
rect 55655 -7369 55707 -7359
rect 55898 -7309 56997 -7308
rect 55898 -7330 56036 -7309
rect 55846 -7370 55898 -7360
rect 56088 -7311 56997 -7309
rect 56088 -7313 56808 -7311
rect 56088 -7330 56230 -7313
rect 56036 -7371 56088 -7361
rect 56282 -7314 56808 -7313
rect 56282 -7315 56616 -7314
rect 56282 -7330 56422 -7315
rect 56230 -7375 56282 -7365
rect 56474 -7330 56616 -7315
rect 56422 -7377 56474 -7367
rect 56668 -7330 56808 -7314
rect 56616 -7376 56668 -7366
rect 56860 -7330 56997 -7311
rect 56808 -7373 56860 -7363
rect 57049 -7330 57191 -7308
rect 56997 -7370 57049 -7360
rect 57243 -7307 66470 -7306
rect 57243 -7330 57384 -7307
rect 57191 -7368 57243 -7358
rect 57436 -7308 58726 -7307
rect 57436 -7330 57577 -7308
rect 57384 -7369 57436 -7359
rect 57629 -7330 57766 -7308
rect 57577 -7370 57629 -7360
rect 57818 -7330 57959 -7308
rect 57766 -7370 57818 -7360
rect 58011 -7330 58151 -7308
rect 57959 -7370 58011 -7360
rect 58203 -7330 58342 -7308
rect 58151 -7370 58203 -7360
rect 58394 -7330 58535 -7308
rect 58342 -7370 58394 -7360
rect 58587 -7330 58726 -7308
rect 58535 -7370 58587 -7360
rect 58778 -7308 61415 -7307
rect 58778 -7330 58921 -7308
rect 58726 -7369 58778 -7359
rect 58973 -7330 59110 -7308
rect 58921 -7370 58973 -7360
rect 59162 -7330 59303 -7308
rect 59110 -7370 59162 -7360
rect 59355 -7330 59495 -7308
rect 59303 -7370 59355 -7360
rect 59547 -7330 59686 -7308
rect 59495 -7370 59547 -7360
rect 59738 -7330 59878 -7308
rect 59686 -7370 59738 -7360
rect 59930 -7330 60071 -7308
rect 59878 -7370 59930 -7360
rect 60123 -7309 60454 -7308
rect 60123 -7330 60260 -7309
rect 60071 -7370 60123 -7360
rect 60312 -7330 60454 -7309
rect 60260 -7371 60312 -7361
rect 60506 -7330 60645 -7308
rect 60454 -7370 60506 -7360
rect 60697 -7330 60838 -7308
rect 60645 -7370 60697 -7360
rect 60890 -7330 61030 -7308
rect 60838 -7370 60890 -7360
rect 61082 -7309 61415 -7308
rect 61082 -7330 61222 -7309
rect 61030 -7370 61082 -7360
rect 61274 -7330 61415 -7309
rect 61222 -7371 61274 -7361
rect 61467 -7330 61605 -7307
rect 61415 -7369 61467 -7359
rect 61657 -7308 62183 -7307
rect 61657 -7309 61990 -7308
rect 61657 -7330 61798 -7309
rect 61605 -7369 61657 -7359
rect 61850 -7330 61990 -7309
rect 61798 -7371 61850 -7361
rect 62042 -7330 62183 -7308
rect 61990 -7370 62042 -7360
rect 62235 -7330 62374 -7307
rect 62183 -7369 62235 -7359
rect 62426 -7308 63143 -7307
rect 62426 -7330 62566 -7308
rect 62374 -7369 62426 -7359
rect 62618 -7330 62757 -7308
rect 62566 -7370 62618 -7360
rect 62809 -7330 62949 -7308
rect 62757 -7370 62809 -7360
rect 63001 -7330 63143 -7308
rect 62949 -7370 63001 -7360
rect 63195 -7308 64102 -7307
rect 63195 -7330 63335 -7308
rect 63143 -7369 63195 -7359
rect 63387 -7309 63909 -7308
rect 63387 -7330 63525 -7309
rect 63335 -7370 63387 -7360
rect 63577 -7310 63909 -7309
rect 63577 -7330 63716 -7310
rect 63525 -7371 63577 -7361
rect 63768 -7330 63909 -7310
rect 63716 -7372 63768 -7362
rect 63961 -7330 64102 -7308
rect 63909 -7370 63961 -7360
rect 64154 -7308 65445 -7307
rect 64154 -7330 64295 -7308
rect 64102 -7369 64154 -7359
rect 64347 -7330 64486 -7308
rect 64295 -7370 64347 -7360
rect 64538 -7330 64677 -7308
rect 64486 -7370 64538 -7360
rect 64729 -7330 64870 -7308
rect 64677 -7370 64729 -7360
rect 64922 -7330 65063 -7308
rect 64870 -7370 64922 -7360
rect 65115 -7330 65254 -7308
rect 65063 -7370 65115 -7360
rect 65306 -7330 65445 -7308
rect 65254 -7370 65306 -7360
rect 65497 -7330 65636 -7307
rect 65445 -7369 65497 -7359
rect 65688 -7308 66470 -7307
rect 65688 -7330 65829 -7308
rect 65636 -7369 65688 -7359
rect 65881 -7330 66023 -7308
rect 65829 -7370 65881 -7360
rect 66075 -7309 66470 -7308
rect 66075 -7330 66211 -7309
rect 66023 -7370 66075 -7360
rect 66263 -7317 66470 -7309
rect 66263 -7330 66405 -7317
rect 66211 -7371 66263 -7361
rect 66457 -7330 66470 -7317
rect 66405 -7379 66457 -7369
rect 49991 -7445 50043 -7435
rect 50182 -7447 50234 -7437
rect 50043 -7490 50182 -7460
rect 50043 -7497 50070 -7490
rect 49991 -7507 50070 -7497
rect 50000 -7654 50070 -7507
rect 50374 -7446 50426 -7436
rect 50234 -7490 50374 -7460
rect 50182 -7509 50234 -7499
rect 50566 -7449 50618 -7439
rect 50426 -7490 50566 -7460
rect 50374 -7508 50426 -7498
rect 50760 -7448 50812 -7438
rect 50618 -7490 50760 -7460
rect 50566 -7511 50618 -7501
rect 50950 -7448 51002 -7438
rect 50812 -7490 50950 -7460
rect 50760 -7510 50812 -7500
rect 51145 -7446 51197 -7436
rect 51002 -7490 51145 -7460
rect 50950 -7510 51002 -7500
rect 51336 -7445 51388 -7435
rect 51197 -7490 51336 -7460
rect 51145 -7508 51197 -7498
rect 51531 -7447 51583 -7437
rect 51388 -7490 51531 -7460
rect 51336 -7507 51388 -7497
rect 51721 -7447 51773 -7437
rect 51583 -7490 51721 -7460
rect 51531 -7509 51583 -7499
rect 51911 -7446 51963 -7436
rect 51773 -7490 51911 -7460
rect 51721 -7509 51773 -7499
rect 52104 -7445 52156 -7435
rect 51963 -7490 52104 -7460
rect 51911 -7508 51963 -7498
rect 52295 -7445 52347 -7435
rect 52156 -7490 52295 -7460
rect 52104 -7507 52156 -7497
rect 52491 -7447 52543 -7437
rect 52347 -7490 52491 -7460
rect 52295 -7507 52347 -7497
rect 52680 -7447 52732 -7437
rect 52543 -7490 52680 -7460
rect 52491 -7509 52543 -7499
rect 52874 -7447 52926 -7437
rect 52732 -7490 52874 -7460
rect 52680 -7509 52732 -7499
rect 53063 -7447 53115 -7437
rect 52926 -7490 53063 -7460
rect 52874 -7509 52926 -7499
rect 53255 -7448 53307 -7438
rect 53115 -7490 53255 -7460
rect 53063 -7509 53115 -7499
rect 53448 -7448 53500 -7438
rect 53307 -7490 53448 -7460
rect 53255 -7510 53307 -7500
rect 53639 -7448 53691 -7438
rect 53500 -7490 53639 -7460
rect 53448 -7510 53500 -7500
rect 53831 -7447 53883 -7437
rect 53691 -7490 53831 -7460
rect 53639 -7510 53691 -7500
rect 54023 -7448 54075 -7438
rect 53883 -7490 54023 -7460
rect 53831 -7509 53883 -7499
rect 54216 -7448 54268 -7438
rect 54075 -7490 54216 -7460
rect 54023 -7510 54075 -7500
rect 54407 -7448 54459 -7438
rect 54268 -7490 54407 -7460
rect 54216 -7510 54268 -7500
rect 54599 -7447 54651 -7437
rect 54459 -7490 54599 -7460
rect 54407 -7510 54459 -7500
rect 54792 -7448 54844 -7438
rect 54651 -7490 54792 -7460
rect 54599 -7509 54651 -7499
rect 54984 -7448 55036 -7438
rect 54844 -7490 54984 -7460
rect 54792 -7510 54844 -7500
rect 55175 -7448 55227 -7438
rect 55036 -7490 55175 -7460
rect 54984 -7510 55036 -7500
rect 55366 -7448 55418 -7438
rect 55227 -7490 55366 -7460
rect 55175 -7510 55227 -7500
rect 55558 -7448 55610 -7438
rect 55418 -7490 55558 -7460
rect 55366 -7510 55418 -7500
rect 55751 -7447 55803 -7437
rect 55610 -7490 55751 -7460
rect 55558 -7510 55610 -7500
rect 55942 -7447 55994 -7437
rect 55803 -7490 55942 -7460
rect 55751 -7509 55803 -7499
rect 56136 -7448 56188 -7438
rect 55994 -7490 56136 -7460
rect 55942 -7509 55994 -7499
rect 56328 -7448 56380 -7438
rect 56188 -7490 56328 -7460
rect 56136 -7510 56188 -7500
rect 56520 -7448 56572 -7438
rect 56380 -7490 56520 -7460
rect 56328 -7510 56380 -7500
rect 56712 -7448 56764 -7438
rect 56572 -7490 56712 -7460
rect 56520 -7510 56572 -7500
rect 56904 -7448 56956 -7438
rect 56764 -7490 56904 -7460
rect 56712 -7510 56764 -7500
rect 57096 -7448 57148 -7438
rect 56956 -7490 57096 -7460
rect 56904 -7510 56956 -7500
rect 57288 -7448 57340 -7438
rect 57148 -7490 57288 -7460
rect 57096 -7510 57148 -7500
rect 57479 -7448 57531 -7438
rect 57340 -7490 57479 -7460
rect 57288 -7510 57340 -7500
rect 57671 -7448 57723 -7438
rect 57531 -7490 57671 -7460
rect 57479 -7510 57531 -7500
rect 57864 -7448 57916 -7438
rect 57723 -7490 57864 -7460
rect 57671 -7510 57723 -7500
rect 58056 -7448 58108 -7438
rect 57916 -7490 58056 -7460
rect 57864 -7510 57916 -7500
rect 58248 -7448 58300 -7438
rect 58108 -7490 58248 -7460
rect 58056 -7510 58108 -7500
rect 58439 -7448 58491 -7438
rect 58300 -7490 58439 -7460
rect 58248 -7510 58300 -7500
rect 58631 -7448 58683 -7438
rect 58491 -7490 58631 -7460
rect 58439 -7510 58491 -7500
rect 58822 -7448 58874 -7438
rect 58683 -7490 58822 -7460
rect 58631 -7510 58683 -7500
rect 59013 -7448 59065 -7438
rect 58874 -7490 59013 -7460
rect 58822 -7510 58874 -7500
rect 59207 -7448 59259 -7438
rect 59065 -7490 59207 -7460
rect 59013 -7510 59065 -7500
rect 59399 -7448 59451 -7438
rect 59259 -7490 59399 -7460
rect 59207 -7510 59259 -7500
rect 59592 -7447 59644 -7437
rect 59451 -7490 59592 -7460
rect 59399 -7510 59451 -7500
rect 59783 -7448 59835 -7438
rect 59644 -7490 59783 -7460
rect 59592 -7509 59644 -7499
rect 59975 -7448 60027 -7438
rect 59835 -7490 59975 -7460
rect 59783 -7510 59835 -7500
rect 60168 -7448 60220 -7438
rect 60027 -7490 60168 -7460
rect 59975 -7510 60027 -7500
rect 60360 -7448 60412 -7438
rect 60220 -7490 60360 -7460
rect 60168 -7510 60220 -7500
rect 60553 -7447 60605 -7437
rect 60412 -7490 60553 -7460
rect 60360 -7510 60412 -7500
rect 60744 -7448 60796 -7438
rect 60605 -7490 60744 -7460
rect 60553 -7509 60605 -7499
rect 60936 -7448 60988 -7438
rect 60796 -7490 60936 -7460
rect 60744 -7510 60796 -7500
rect 61127 -7448 61179 -7438
rect 60988 -7490 61127 -7460
rect 60936 -7510 60988 -7500
rect 61319 -7448 61371 -7438
rect 61179 -7490 61319 -7460
rect 61127 -7510 61179 -7500
rect 61511 -7448 61563 -7438
rect 61371 -7490 61511 -7460
rect 61319 -7510 61371 -7500
rect 61704 -7448 61756 -7438
rect 61563 -7490 61704 -7460
rect 61511 -7510 61563 -7500
rect 61895 -7448 61947 -7438
rect 61756 -7490 61895 -7460
rect 61704 -7510 61756 -7500
rect 62087 -7448 62139 -7438
rect 61947 -7490 62087 -7460
rect 61895 -7510 61947 -7500
rect 62279 -7447 62331 -7437
rect 62139 -7490 62279 -7460
rect 62087 -7510 62139 -7500
rect 62471 -7448 62523 -7438
rect 62331 -7490 62471 -7460
rect 62279 -7509 62331 -7499
rect 62661 -7448 62713 -7438
rect 62523 -7490 62661 -7460
rect 62471 -7510 62523 -7500
rect 62855 -7448 62907 -7438
rect 62713 -7490 62855 -7460
rect 62661 -7510 62713 -7500
rect 63047 -7447 63099 -7437
rect 62907 -7490 63047 -7460
rect 62855 -7510 62907 -7500
rect 63238 -7448 63290 -7438
rect 63099 -7490 63238 -7460
rect 63047 -7509 63099 -7499
rect 63431 -7448 63483 -7438
rect 63290 -7490 63431 -7460
rect 63238 -7510 63290 -7500
rect 63622 -7447 63674 -7437
rect 63483 -7490 63622 -7460
rect 63431 -7510 63483 -7500
rect 63814 -7448 63866 -7438
rect 63674 -7490 63814 -7460
rect 63622 -7509 63674 -7499
rect 64005 -7448 64057 -7438
rect 63866 -7490 64005 -7460
rect 63814 -7510 63866 -7500
rect 64199 -7447 64251 -7437
rect 64057 -7490 64199 -7460
rect 64005 -7510 64057 -7500
rect 64390 -7448 64442 -7438
rect 64251 -7490 64390 -7460
rect 64199 -7509 64251 -7499
rect 64582 -7448 64634 -7438
rect 64442 -7490 64582 -7460
rect 64390 -7510 64442 -7500
rect 64774 -7448 64826 -7438
rect 64634 -7490 64774 -7460
rect 64582 -7510 64634 -7500
rect 64966 -7448 65018 -7438
rect 64826 -7490 64966 -7460
rect 64774 -7510 64826 -7500
rect 65159 -7448 65211 -7438
rect 65018 -7490 65159 -7460
rect 64966 -7510 65018 -7500
rect 65350 -7448 65402 -7438
rect 65211 -7490 65350 -7460
rect 65159 -7510 65211 -7500
rect 65543 -7447 65595 -7437
rect 65402 -7490 65543 -7460
rect 65350 -7510 65402 -7500
rect 65734 -7448 65786 -7438
rect 65595 -7490 65734 -7460
rect 65543 -7509 65595 -7499
rect 65927 -7448 65979 -7438
rect 65786 -7490 65927 -7460
rect 65734 -7510 65786 -7500
rect 66118 -7448 66170 -7438
rect 65979 -7490 66118 -7460
rect 65927 -7510 65979 -7500
rect 66309 -7446 66361 -7436
rect 66170 -7490 66309 -7460
rect 66118 -7510 66170 -7500
rect 66504 -7448 66556 -7438
rect 66361 -7490 66504 -7460
rect 66309 -7508 66361 -7498
rect 66440 -7500 66504 -7490
rect 66440 -7510 66556 -7500
rect 66440 -7654 66510 -7510
rect 49940 -7664 66588 -7654
rect 47224 -7808 47652 -7752
rect 48274 -7706 48446 -7696
rect 48274 -7774 48446 -7764
rect 49940 -7766 66588 -7756
rect 68120 -7710 68292 -7700
rect 68120 -7778 68292 -7768
rect 68894 -7756 68924 -6672
rect 69290 -7756 69326 -6672
rect 68894 -7806 69326 -7756
rect 68584 -7808 69326 -7806
rect 47224 -8196 69326 -7808
rect 47482 -8198 69326 -8196
<< via2 >>
rect 48286 -5236 48444 -5178
rect 49920 -5280 66554 -5188
rect 68070 -5236 68228 -5178
rect 51516 -6364 51572 -6308
rect 51720 -6618 51776 -6562
rect 51938 -6354 51994 -6298
rect 52330 -6354 52386 -6298
rect 52716 -6342 52772 -6286
rect 53102 -6344 53158 -6288
rect 52132 -6490 52188 -6434
rect 52510 -6488 52566 -6432
rect 53486 -6352 53542 -6296
rect 53872 -6350 53928 -6294
rect 52908 -6488 52964 -6432
rect 53294 -6490 53350 -6434
rect 54256 -6352 54312 -6296
rect 54638 -6354 54694 -6298
rect 55018 -6348 55074 -6292
rect 55412 -6360 55468 -6304
rect 55782 -6358 55838 -6302
rect 53672 -6490 53728 -6434
rect 54056 -6492 54112 -6436
rect 54428 -6492 54484 -6436
rect 54820 -6492 54876 -6436
rect 55198 -6492 55254 -6436
rect 56174 -6354 56230 -6298
rect 55594 -6488 55650 -6432
rect 56560 -6356 56616 -6300
rect 56936 -6352 56992 -6296
rect 57312 -6356 57368 -6300
rect 57708 -6354 57764 -6298
rect 58128 -6348 58184 -6292
rect 58520 -6350 58576 -6294
rect 58908 -6350 58964 -6294
rect 59290 -6354 59346 -6298
rect 55974 -6490 56030 -6434
rect 56352 -6492 56408 -6436
rect 56744 -6492 56800 -6436
rect 57126 -6492 57182 -6436
rect 57500 -6492 57556 -6436
rect 58322 -6492 58378 -6436
rect 58712 -6492 58768 -6436
rect 59690 -6352 59746 -6296
rect 60066 -6346 60122 -6290
rect 60438 -6350 60494 -6294
rect 60836 -6356 60892 -6300
rect 61218 -6352 61274 -6296
rect 61592 -6350 61648 -6294
rect 59100 -6490 59156 -6434
rect 59490 -6492 59546 -6436
rect 59858 -6492 59914 -6436
rect 60252 -6492 60308 -6436
rect 60644 -6490 60700 -6434
rect 61010 -6490 61066 -6434
rect 61972 -6352 62028 -6296
rect 62360 -6352 62416 -6296
rect 61406 -6488 61462 -6432
rect 61782 -6492 61838 -6436
rect 62742 -6350 62798 -6294
rect 63128 -6352 63184 -6296
rect 62162 -6490 62218 -6434
rect 62550 -6492 62606 -6436
rect 63510 -6350 63566 -6294
rect 63898 -6348 63954 -6292
rect 62936 -6490 62992 -6434
rect 63316 -6492 63372 -6436
rect 63706 -6490 63762 -6434
rect 52238 -6618 52294 -6562
rect 51838 -6746 51894 -6690
rect 52044 -6746 52100 -6690
rect 52620 -6618 52676 -6562
rect 52432 -6752 52488 -6696
rect 53002 -6618 53058 -6562
rect 52818 -6748 52874 -6692
rect 53390 -6618 53446 -6562
rect 53200 -6746 53256 -6690
rect 53768 -6618 53824 -6562
rect 53582 -6748 53638 -6692
rect 54150 -6618 54206 -6562
rect 53964 -6750 54020 -6694
rect 54538 -6618 54594 -6562
rect 54350 -6750 54406 -6694
rect 54920 -6618 54976 -6562
rect 54740 -6748 54796 -6692
rect 55304 -6618 55360 -6562
rect 55120 -6752 55176 -6696
rect 55682 -6618 55738 -6562
rect 56072 -6618 56128 -6562
rect 55502 -6752 55558 -6696
rect 55886 -6750 55942 -6694
rect 56454 -6618 56510 -6562
rect 56272 -6748 56328 -6692
rect 56840 -6618 56896 -6562
rect 57222 -6618 57278 -6562
rect 56658 -6750 56714 -6694
rect 57038 -6752 57094 -6696
rect 57602 -6618 57658 -6562
rect 57422 -6752 57478 -6696
rect 58414 -6618 58470 -6562
rect 58796 -6618 58852 -6562
rect 57806 -6750 57862 -6694
rect 58230 -6750 58286 -6694
rect 58612 -6754 58668 -6698
rect 59186 -6618 59242 -6562
rect 58996 -6750 59052 -6694
rect 59568 -6618 59624 -6562
rect 59382 -6750 59438 -6694
rect 59954 -6618 60010 -6562
rect 59764 -6750 59820 -6694
rect 60336 -6618 60392 -6562
rect 60154 -6748 60210 -6692
rect 60722 -6618 60778 -6562
rect 60534 -6752 60590 -6696
rect 61104 -6618 61160 -6562
rect 60918 -6750 60974 -6694
rect 61482 -6618 61538 -6562
rect 61866 -6618 61922 -6562
rect 62252 -6618 62308 -6562
rect 62640 -6618 62696 -6562
rect 61300 -6750 61356 -6694
rect 61688 -6752 61744 -6696
rect 62070 -6748 62126 -6692
rect 62456 -6748 62512 -6692
rect 63022 -6618 63078 -6562
rect 62840 -6746 62896 -6690
rect 63406 -6618 63462 -6562
rect 63220 -6748 63276 -6692
rect 63792 -6618 63848 -6562
rect 63608 -6746 63664 -6690
rect 64502 -6492 64558 -6436
rect 64238 -6618 64294 -6562
rect 63992 -6746 64048 -6690
rect 64144 -6746 64200 -6690
rect 48274 -7764 48432 -7706
rect 49940 -7756 66574 -7664
rect 68120 -7768 68278 -7710
<< metal3 >>
rect 62104 -5160 62384 -5150
rect 67454 -5160 67734 -5150
rect 46340 -5178 69982 -5160
rect 46340 -5236 48286 -5178
rect 48444 -5188 68070 -5178
rect 48444 -5236 49920 -5188
rect 46340 -5280 49920 -5236
rect 66554 -5236 68070 -5188
rect 68228 -5236 69982 -5178
rect 66554 -5280 69982 -5236
rect 46340 -5438 69982 -5280
rect 52706 -6286 52782 -6281
rect 51928 -6298 52004 -6293
rect 51506 -6304 51582 -6303
rect 51928 -6304 51938 -6298
rect 51506 -6308 51938 -6304
rect 51506 -6364 51516 -6308
rect 51572 -6354 51938 -6308
rect 51994 -6304 52004 -6298
rect 52320 -6298 52396 -6293
rect 52320 -6304 52330 -6298
rect 51994 -6354 52330 -6304
rect 52386 -6304 52396 -6298
rect 52706 -6304 52716 -6286
rect 52386 -6342 52716 -6304
rect 52772 -6304 52782 -6286
rect 53092 -6288 53168 -6283
rect 53092 -6304 53102 -6288
rect 52772 -6342 53102 -6304
rect 52386 -6344 53102 -6342
rect 53158 -6304 53168 -6288
rect 53476 -6296 53552 -6291
rect 53476 -6304 53486 -6296
rect 53158 -6344 53486 -6304
rect 52386 -6352 53486 -6344
rect 53542 -6304 53552 -6296
rect 53862 -6294 53938 -6289
rect 53862 -6304 53872 -6294
rect 53542 -6350 53872 -6304
rect 53928 -6304 53938 -6294
rect 54246 -6296 54322 -6291
rect 55008 -6292 55084 -6287
rect 54246 -6304 54256 -6296
rect 53928 -6350 54256 -6304
rect 53542 -6352 54256 -6350
rect 54312 -6304 54322 -6296
rect 54628 -6298 54704 -6293
rect 54628 -6304 54638 -6298
rect 54312 -6352 54638 -6304
rect 52386 -6354 54638 -6352
rect 54694 -6304 54704 -6298
rect 55008 -6304 55018 -6292
rect 54694 -6348 55018 -6304
rect 55074 -6304 55084 -6292
rect 55402 -6304 55478 -6299
rect 55772 -6302 55848 -6297
rect 55772 -6304 55782 -6302
rect 55074 -6348 55412 -6304
rect 54694 -6354 55412 -6348
rect 51572 -6360 55412 -6354
rect 55468 -6358 55782 -6304
rect 55838 -6304 55848 -6302
rect 56164 -6298 56240 -6293
rect 56164 -6304 56174 -6298
rect 55838 -6354 56174 -6304
rect 56230 -6304 56240 -6298
rect 56550 -6300 56626 -6295
rect 56550 -6304 56560 -6300
rect 56230 -6354 56560 -6304
rect 55838 -6356 56560 -6354
rect 56616 -6304 56626 -6300
rect 56926 -6296 57002 -6291
rect 58118 -6292 58194 -6287
rect 56926 -6304 56936 -6296
rect 56616 -6352 56936 -6304
rect 56992 -6304 57002 -6296
rect 57302 -6300 57378 -6295
rect 57302 -6304 57312 -6300
rect 56992 -6352 57312 -6304
rect 56616 -6356 57312 -6352
rect 57368 -6304 57378 -6300
rect 57698 -6298 57774 -6293
rect 57698 -6304 57708 -6298
rect 57368 -6354 57708 -6304
rect 57764 -6304 57774 -6298
rect 58118 -6304 58128 -6292
rect 57764 -6348 58128 -6304
rect 58184 -6304 58194 -6292
rect 58510 -6294 58586 -6289
rect 58510 -6304 58520 -6294
rect 58184 -6348 58520 -6304
rect 57764 -6350 58520 -6348
rect 58576 -6304 58586 -6294
rect 58898 -6294 58974 -6289
rect 60056 -6290 60132 -6285
rect 58898 -6304 58908 -6294
rect 58576 -6350 58908 -6304
rect 58964 -6304 58974 -6294
rect 59280 -6298 59356 -6293
rect 59280 -6304 59290 -6298
rect 58964 -6350 59290 -6304
rect 57764 -6354 59290 -6350
rect 59346 -6304 59356 -6298
rect 59680 -6296 59756 -6291
rect 59680 -6304 59690 -6296
rect 59346 -6352 59690 -6304
rect 59746 -6304 59756 -6296
rect 60056 -6304 60066 -6290
rect 59746 -6346 60066 -6304
rect 60122 -6304 60132 -6290
rect 60428 -6294 60504 -6289
rect 60428 -6304 60438 -6294
rect 60122 -6346 60438 -6304
rect 59746 -6350 60438 -6346
rect 60494 -6304 60504 -6294
rect 60826 -6300 60902 -6295
rect 60826 -6304 60836 -6300
rect 60494 -6350 60836 -6304
rect 59746 -6352 60836 -6350
rect 59346 -6354 60836 -6352
rect 57368 -6356 60836 -6354
rect 60892 -6304 60902 -6300
rect 61208 -6296 61284 -6291
rect 61208 -6304 61218 -6296
rect 60892 -6352 61218 -6304
rect 61274 -6304 61284 -6296
rect 61582 -6294 61658 -6289
rect 61582 -6304 61592 -6294
rect 61274 -6350 61592 -6304
rect 61648 -6304 61658 -6294
rect 61962 -6296 62038 -6291
rect 61962 -6304 61972 -6296
rect 61648 -6350 61972 -6304
rect 61274 -6352 61972 -6350
rect 62028 -6304 62038 -6296
rect 62350 -6296 62426 -6291
rect 62350 -6304 62360 -6296
rect 62028 -6352 62360 -6304
rect 62416 -6304 62426 -6296
rect 62732 -6294 62808 -6289
rect 62732 -6304 62742 -6294
rect 62416 -6350 62742 -6304
rect 62798 -6304 62808 -6294
rect 63118 -6296 63194 -6291
rect 63118 -6304 63128 -6296
rect 62798 -6350 63128 -6304
rect 62416 -6352 63128 -6350
rect 63184 -6304 63194 -6296
rect 63500 -6294 63576 -6289
rect 63500 -6304 63510 -6294
rect 63184 -6350 63510 -6304
rect 63566 -6304 63576 -6294
rect 63888 -6292 63964 -6287
rect 63888 -6304 63898 -6292
rect 63566 -6348 63898 -6304
rect 63954 -6304 63964 -6292
rect 63954 -6348 64124 -6304
rect 63566 -6350 64124 -6348
rect 63184 -6352 64124 -6350
rect 60892 -6356 64124 -6352
rect 55838 -6358 64124 -6356
rect 55468 -6360 64124 -6358
rect 51572 -6364 64124 -6360
rect 51506 -6366 64124 -6364
rect 51506 -6369 51582 -6366
rect 52122 -6434 52198 -6429
rect 52500 -6432 52576 -6427
rect 52500 -6434 52510 -6432
rect 51918 -6490 52132 -6434
rect 52188 -6488 52510 -6434
rect 52566 -6434 52576 -6432
rect 52898 -6432 52974 -6427
rect 52898 -6434 52908 -6432
rect 52566 -6488 52908 -6434
rect 52964 -6434 52974 -6432
rect 53284 -6434 53360 -6429
rect 53662 -6434 53738 -6429
rect 54046 -6434 54122 -6431
rect 54418 -6434 54494 -6431
rect 54810 -6434 54886 -6431
rect 55188 -6434 55264 -6431
rect 55584 -6432 55660 -6427
rect 55584 -6434 55594 -6432
rect 52964 -6488 53294 -6434
rect 52188 -6490 53294 -6488
rect 53350 -6490 53672 -6434
rect 53728 -6436 55594 -6434
rect 53728 -6490 54056 -6436
rect 51918 -6492 54056 -6490
rect 54112 -6492 54428 -6436
rect 54484 -6492 54820 -6436
rect 54876 -6492 55198 -6436
rect 55254 -6488 55594 -6436
rect 55650 -6434 55660 -6432
rect 55964 -6434 56040 -6429
rect 56342 -6434 56418 -6431
rect 56734 -6434 56810 -6431
rect 57116 -6434 57192 -6431
rect 57490 -6434 57566 -6431
rect 58312 -6434 58388 -6431
rect 58702 -6434 58778 -6431
rect 59090 -6434 59166 -6429
rect 59480 -6434 59556 -6431
rect 59848 -6434 59924 -6431
rect 60242 -6434 60318 -6431
rect 60634 -6434 60710 -6429
rect 61000 -6434 61076 -6429
rect 61396 -6432 61472 -6427
rect 61396 -6434 61406 -6432
rect 55650 -6488 55974 -6434
rect 55254 -6490 55974 -6488
rect 56030 -6436 59100 -6434
rect 56030 -6490 56352 -6436
rect 55254 -6492 56352 -6490
rect 56408 -6492 56744 -6436
rect 56800 -6492 57126 -6436
rect 57182 -6492 57500 -6436
rect 57556 -6492 58322 -6436
rect 58378 -6492 58712 -6436
rect 58768 -6490 59100 -6436
rect 59156 -6436 60644 -6434
rect 59156 -6490 59490 -6436
rect 58768 -6492 59490 -6490
rect 59546 -6492 59858 -6436
rect 59914 -6492 60252 -6436
rect 60308 -6490 60644 -6436
rect 60700 -6490 61010 -6434
rect 61066 -6488 61406 -6434
rect 61462 -6434 61472 -6432
rect 61772 -6434 61848 -6431
rect 62152 -6434 62228 -6429
rect 62540 -6434 62616 -6431
rect 62926 -6434 63002 -6429
rect 63306 -6434 63382 -6431
rect 63696 -6434 63772 -6429
rect 64492 -6434 64568 -6431
rect 61462 -6436 62162 -6434
rect 61462 -6488 61782 -6436
rect 61066 -6490 61782 -6488
rect 60308 -6492 61782 -6490
rect 61838 -6490 62162 -6436
rect 62218 -6436 62936 -6434
rect 62218 -6490 62550 -6436
rect 61838 -6492 62550 -6490
rect 62606 -6490 62936 -6436
rect 62992 -6436 63706 -6434
rect 62992 -6490 63316 -6436
rect 62606 -6492 63316 -6490
rect 63372 -6490 63706 -6436
rect 63762 -6436 64568 -6434
rect 63762 -6490 64502 -6436
rect 63372 -6492 64502 -6490
rect 64558 -6492 64568 -6436
rect 51918 -6496 64568 -6492
rect 54046 -6497 54122 -6496
rect 54418 -6497 54494 -6496
rect 54810 -6497 54886 -6496
rect 55188 -6497 55264 -6496
rect 56342 -6497 56418 -6496
rect 56734 -6497 56810 -6496
rect 57116 -6497 57192 -6496
rect 57490 -6497 57566 -6496
rect 58312 -6497 58388 -6496
rect 58702 -6497 58778 -6496
rect 59480 -6497 59556 -6496
rect 59848 -6497 59924 -6496
rect 60242 -6497 60318 -6496
rect 61772 -6497 61848 -6496
rect 62540 -6497 62616 -6496
rect 63306 -6497 63382 -6496
rect 64492 -6497 64568 -6496
rect 51710 -6562 51786 -6557
rect 52228 -6562 52304 -6557
rect 52610 -6562 52686 -6557
rect 52992 -6562 53068 -6557
rect 53380 -6562 53456 -6557
rect 53758 -6562 53834 -6557
rect 54140 -6562 54216 -6557
rect 54528 -6562 54604 -6557
rect 54910 -6562 54986 -6557
rect 55294 -6562 55370 -6557
rect 55672 -6562 55748 -6557
rect 56062 -6562 56138 -6557
rect 56444 -6562 56520 -6557
rect 56830 -6562 56906 -6557
rect 57212 -6562 57288 -6557
rect 57592 -6562 57668 -6557
rect 58404 -6562 58480 -6557
rect 58786 -6562 58862 -6557
rect 59176 -6562 59252 -6557
rect 59558 -6562 59634 -6557
rect 59944 -6562 60020 -6557
rect 60326 -6562 60402 -6557
rect 60712 -6562 60788 -6557
rect 61094 -6562 61170 -6557
rect 61472 -6562 61548 -6557
rect 61856 -6562 61932 -6557
rect 62242 -6562 62318 -6557
rect 62630 -6562 62706 -6557
rect 63012 -6562 63088 -6557
rect 63396 -6562 63472 -6557
rect 63782 -6562 63858 -6557
rect 64228 -6562 64304 -6557
rect 51692 -6618 51720 -6562
rect 51776 -6618 52238 -6562
rect 52294 -6618 52620 -6562
rect 52676 -6618 53002 -6562
rect 53058 -6618 53390 -6562
rect 53446 -6618 53768 -6562
rect 53824 -6618 54150 -6562
rect 54206 -6618 54538 -6562
rect 54594 -6618 54920 -6562
rect 54976 -6618 55304 -6562
rect 55360 -6618 55682 -6562
rect 55738 -6618 56072 -6562
rect 56128 -6618 56454 -6562
rect 56510 -6618 56840 -6562
rect 56896 -6618 57222 -6562
rect 57278 -6618 57602 -6562
rect 57658 -6618 58414 -6562
rect 58470 -6618 58796 -6562
rect 58852 -6618 59186 -6562
rect 59242 -6618 59568 -6562
rect 59624 -6618 59954 -6562
rect 60010 -6618 60336 -6562
rect 60392 -6618 60722 -6562
rect 60778 -6618 61104 -6562
rect 61160 -6618 61482 -6562
rect 61538 -6618 61866 -6562
rect 61922 -6618 62252 -6562
rect 62308 -6618 62640 -6562
rect 62696 -6618 63022 -6562
rect 63078 -6618 63406 -6562
rect 63462 -6618 63792 -6562
rect 63848 -6618 64238 -6562
rect 64294 -6618 64332 -6562
rect 51692 -6624 64332 -6618
rect 51684 -6690 64330 -6684
rect 51684 -6746 51838 -6690
rect 51894 -6746 52044 -6690
rect 52100 -6692 53200 -6690
rect 52100 -6696 52818 -6692
rect 52100 -6746 52432 -6696
rect 51828 -6751 51904 -6746
rect 52034 -6751 52110 -6746
rect 52422 -6752 52432 -6746
rect 52488 -6746 52818 -6696
rect 52488 -6752 52498 -6746
rect 52422 -6757 52498 -6752
rect 52808 -6748 52818 -6746
rect 52874 -6746 53200 -6692
rect 53256 -6692 62840 -6690
rect 53256 -6746 53582 -6692
rect 52874 -6748 52884 -6746
rect 52808 -6753 52884 -6748
rect 53190 -6751 53266 -6746
rect 53572 -6748 53582 -6746
rect 53638 -6694 54740 -6692
rect 53638 -6746 53964 -6694
rect 53638 -6748 53648 -6746
rect 53572 -6753 53648 -6748
rect 53954 -6750 53964 -6746
rect 54020 -6746 54350 -6694
rect 54020 -6750 54030 -6746
rect 53954 -6755 54030 -6750
rect 54340 -6750 54350 -6746
rect 54406 -6746 54740 -6694
rect 54406 -6750 54416 -6746
rect 54340 -6755 54416 -6750
rect 54730 -6748 54740 -6746
rect 54796 -6694 56272 -6692
rect 54796 -6696 55886 -6694
rect 54796 -6746 55120 -6696
rect 54796 -6748 54806 -6746
rect 54730 -6753 54806 -6748
rect 55110 -6752 55120 -6746
rect 55176 -6746 55502 -6696
rect 55176 -6752 55186 -6746
rect 55110 -6757 55186 -6752
rect 55492 -6752 55502 -6746
rect 55558 -6746 55886 -6696
rect 55558 -6752 55568 -6746
rect 55492 -6757 55568 -6752
rect 55876 -6750 55886 -6746
rect 55942 -6746 56272 -6694
rect 55942 -6750 55952 -6746
rect 55876 -6755 55952 -6750
rect 56262 -6748 56272 -6746
rect 56328 -6694 60154 -6692
rect 56328 -6746 56658 -6694
rect 56328 -6748 56338 -6746
rect 56262 -6753 56338 -6748
rect 56648 -6750 56658 -6746
rect 56714 -6696 57806 -6694
rect 56714 -6746 57038 -6696
rect 56714 -6750 56724 -6746
rect 56648 -6755 56724 -6750
rect 57028 -6752 57038 -6746
rect 57094 -6746 57422 -6696
rect 57094 -6752 57104 -6746
rect 57028 -6757 57104 -6752
rect 57412 -6752 57422 -6746
rect 57478 -6746 57806 -6696
rect 57478 -6752 57488 -6746
rect 57412 -6757 57488 -6752
rect 57796 -6750 57806 -6746
rect 57862 -6746 58230 -6694
rect 57862 -6750 57872 -6746
rect 57796 -6755 57872 -6750
rect 58220 -6750 58230 -6746
rect 58286 -6698 58996 -6694
rect 58286 -6746 58612 -6698
rect 58286 -6750 58296 -6746
rect 58220 -6755 58296 -6750
rect 58602 -6754 58612 -6746
rect 58668 -6746 58996 -6698
rect 58668 -6754 58678 -6746
rect 58602 -6759 58678 -6754
rect 58986 -6750 58996 -6746
rect 59052 -6746 59382 -6694
rect 59052 -6750 59062 -6746
rect 58986 -6755 59062 -6750
rect 59372 -6750 59382 -6746
rect 59438 -6746 59764 -6694
rect 59438 -6750 59448 -6746
rect 59372 -6755 59448 -6750
rect 59754 -6750 59764 -6746
rect 59820 -6746 60154 -6694
rect 59820 -6750 59830 -6746
rect 59754 -6755 59830 -6750
rect 60144 -6748 60154 -6746
rect 60210 -6694 62070 -6692
rect 60210 -6696 60918 -6694
rect 60210 -6746 60534 -6696
rect 60210 -6748 60220 -6746
rect 60144 -6753 60220 -6748
rect 60524 -6752 60534 -6746
rect 60590 -6746 60918 -6696
rect 60590 -6752 60600 -6746
rect 60524 -6757 60600 -6752
rect 60908 -6750 60918 -6746
rect 60974 -6746 61300 -6694
rect 60974 -6750 60984 -6746
rect 60908 -6755 60984 -6750
rect 61290 -6750 61300 -6746
rect 61356 -6696 62070 -6694
rect 61356 -6746 61688 -6696
rect 61356 -6750 61366 -6746
rect 61290 -6755 61366 -6750
rect 61678 -6752 61688 -6746
rect 61744 -6746 62070 -6696
rect 61744 -6752 61754 -6746
rect 61678 -6757 61754 -6752
rect 62060 -6748 62070 -6746
rect 62126 -6746 62456 -6692
rect 62126 -6748 62136 -6746
rect 62060 -6753 62136 -6748
rect 62446 -6748 62456 -6746
rect 62512 -6746 62840 -6692
rect 62896 -6692 63608 -6690
rect 62896 -6746 63220 -6692
rect 62512 -6748 62522 -6746
rect 62446 -6753 62522 -6748
rect 62830 -6751 62906 -6746
rect 63210 -6748 63220 -6746
rect 63276 -6746 63608 -6692
rect 63664 -6746 63992 -6690
rect 64048 -6746 64144 -6690
rect 64200 -6746 64330 -6690
rect 63276 -6748 63286 -6746
rect 63210 -6753 63286 -6748
rect 63598 -6751 63674 -6746
rect 63982 -6751 64058 -6746
rect 64134 -6751 64210 -6746
rect 46350 -7664 69992 -7510
rect 46350 -7706 49940 -7664
rect 46350 -7764 48274 -7706
rect 48432 -7756 49940 -7706
rect 66574 -7710 69992 -7664
rect 66574 -7756 68120 -7710
rect 48432 -7764 68120 -7756
rect 46350 -7768 68120 -7764
rect 68278 -7768 69992 -7710
rect 46350 -7788 69992 -7768
use sky130_fd_pr__nfet_01v8_lvt_MNZFGM  XM20
timestamp 1672437577
transform 1 0 54907 0 1 -6788
box -2957 -188 2957 188
use sky130_fd_pr__nfet_01v8_lvt_MNZFGM  XM21
timestamp 1672437577
transform 1 0 54901 0 1 -6166
box -2957 -188 2957 188
use sky130_fd_pr__nfet_01v8_lvt_MNZFGM  XM23
timestamp 1672437577
transform 1 0 61089 0 1 -6776
box -2957 -188 2957 188
use sky130_fd_pr__nfet_01v8_lvt_G3ZQK6  XM24
timestamp 1662412052
transform 1 0 58273 0 1 -5540
box -8423 -310 8423 310
use sky130_fd_pr__nfet_01v8_lvt_G3ZQK6  XM25
timestamp 1662412052
transform 1 0 58273 0 1 -7398
box -8423 -310 8423 310
use sky130_fd_pr__res_xhigh_po_5p73_4C7XCD  XR19
timestamp 1662952458
transform 0 1 47715 -1 0 -7211
box -739 -657 739 657
use sky130_fd_pr__res_xhigh_po_5p73_4C7XCD  XR20
timestamp 1662952458
transform 0 1 47715 -1 0 -5727
box -739 -657 739 657
use sky130_fd_pr__res_xhigh_po_5p73_QP6N54  XR21
timestamp 1662952458
transform 1 0 49111 0 1 -6518
box -739 -748 739 748
use sky130_fd_pr__res_xhigh_po_5p73_4C7XCD  XR22
timestamp 1662952458
transform 0 1 68837 -1 0 -5731
box -739 -657 739 657
use sky130_fd_pr__nfet_01v8_lvt_MNZFGM  sky130_fd_pr__nfet_01v8_lvt_MNZFGM_0
timestamp 1672437577
transform 1 0 61095 0 1 -6166
box -2957 -188 2957 188
use sky130_fd_pr__res_xhigh_po_5p73_4C7XCD  sky130_fd_pr__res_xhigh_po_5p73_4C7XCD_0
timestamp 1662952458
transform 0 1 68837 -1 0 -7211
box -739 -657 739 657
use sky130_fd_pr__res_xhigh_po_5p73_QP6N54  sky130_fd_pr__res_xhigh_po_5p73_QP6N54_0
timestamp 1662952458
transform 1 0 67439 0 1 -6468
box -739 -748 739 748
<< labels >>
rlabel metal1 49890 -7550 49890 -7550 7 vc1
port 7 w
rlabel metal1 49880 -5390 49880 -5390 7 vc2
port 8 w
<< end >>
