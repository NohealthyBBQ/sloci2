magic
tech sky130A
magscale 1 2
timestamp 1672530722
<< metal3 >>
rect -120 680 120 737
rect -120 -737 120 -680
<< rmetal3 >>
rect -120 -680 120 680
<< properties >>
string gencell sky130_fd_pr__res_generic_m3
string library sky130
string parameters w 1.2 l 6.8 m 1 nx 1 wmin 0.30 lmin 0.30 rho 0.047 val 266.333m dummy 0 dw 0.0 term 0.0 roverlap 0
<< end >>
