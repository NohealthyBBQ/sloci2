magic
tech sky130A
magscale 1 2
timestamp 1662988209
<< error_p >>
rect -29 2053 29 2059
rect -29 2019 -17 2053
rect -29 2013 29 2019
rect -29 1743 29 1749
rect -29 1709 -17 1743
rect -29 1703 29 1709
rect -29 1635 29 1641
rect -29 1601 -17 1635
rect -29 1595 29 1601
rect -29 1325 29 1331
rect -29 1291 -17 1325
rect -29 1285 29 1291
rect -29 1217 29 1223
rect -29 1183 -17 1217
rect -29 1177 29 1183
rect -29 907 29 913
rect -29 873 -17 907
rect -29 867 29 873
rect -29 799 29 805
rect -29 765 -17 799
rect -29 759 29 765
rect -29 489 29 495
rect -29 455 -17 489
rect -29 449 29 455
rect -29 381 29 387
rect -29 347 -17 381
rect -29 341 29 347
rect -29 71 29 77
rect -29 37 -17 71
rect -29 31 29 37
rect -29 -37 29 -31
rect -29 -71 -17 -37
rect -29 -77 29 -71
rect -29 -347 29 -341
rect -29 -381 -17 -347
rect -29 -387 29 -381
rect -29 -455 29 -449
rect -29 -489 -17 -455
rect -29 -495 29 -489
rect -29 -765 29 -759
rect -29 -799 -17 -765
rect -29 -805 29 -799
rect -29 -873 29 -867
rect -29 -907 -17 -873
rect -29 -913 29 -907
rect -29 -1183 29 -1177
rect -29 -1217 -17 -1183
rect -29 -1223 29 -1217
rect -29 -1291 29 -1285
rect -29 -1325 -17 -1291
rect -29 -1331 29 -1325
rect -29 -1601 29 -1595
rect -29 -1635 -17 -1601
rect -29 -1641 29 -1635
rect -29 -1709 29 -1703
rect -29 -1743 -17 -1709
rect -29 -1749 29 -1743
rect -29 -2019 29 -2013
rect -29 -2053 -17 -2019
rect -29 -2059 29 -2053
<< pwell >>
rect -211 -2191 211 2191
<< nmoslvt >>
rect -15 1781 15 1981
rect -15 1363 15 1563
rect -15 945 15 1145
rect -15 527 15 727
rect -15 109 15 309
rect -15 -309 15 -109
rect -15 -727 15 -527
rect -15 -1145 15 -945
rect -15 -1563 15 -1363
rect -15 -1981 15 -1781
<< ndiff >>
rect -73 1969 -15 1981
rect -73 1793 -61 1969
rect -27 1793 -15 1969
rect -73 1781 -15 1793
rect 15 1969 73 1981
rect 15 1793 27 1969
rect 61 1793 73 1969
rect 15 1781 73 1793
rect -73 1551 -15 1563
rect -73 1375 -61 1551
rect -27 1375 -15 1551
rect -73 1363 -15 1375
rect 15 1551 73 1563
rect 15 1375 27 1551
rect 61 1375 73 1551
rect 15 1363 73 1375
rect -73 1133 -15 1145
rect -73 957 -61 1133
rect -27 957 -15 1133
rect -73 945 -15 957
rect 15 1133 73 1145
rect 15 957 27 1133
rect 61 957 73 1133
rect 15 945 73 957
rect -73 715 -15 727
rect -73 539 -61 715
rect -27 539 -15 715
rect -73 527 -15 539
rect 15 715 73 727
rect 15 539 27 715
rect 61 539 73 715
rect 15 527 73 539
rect -73 297 -15 309
rect -73 121 -61 297
rect -27 121 -15 297
rect -73 109 -15 121
rect 15 297 73 309
rect 15 121 27 297
rect 61 121 73 297
rect 15 109 73 121
rect -73 -121 -15 -109
rect -73 -297 -61 -121
rect -27 -297 -15 -121
rect -73 -309 -15 -297
rect 15 -121 73 -109
rect 15 -297 27 -121
rect 61 -297 73 -121
rect 15 -309 73 -297
rect -73 -539 -15 -527
rect -73 -715 -61 -539
rect -27 -715 -15 -539
rect -73 -727 -15 -715
rect 15 -539 73 -527
rect 15 -715 27 -539
rect 61 -715 73 -539
rect 15 -727 73 -715
rect -73 -957 -15 -945
rect -73 -1133 -61 -957
rect -27 -1133 -15 -957
rect -73 -1145 -15 -1133
rect 15 -957 73 -945
rect 15 -1133 27 -957
rect 61 -1133 73 -957
rect 15 -1145 73 -1133
rect -73 -1375 -15 -1363
rect -73 -1551 -61 -1375
rect -27 -1551 -15 -1375
rect -73 -1563 -15 -1551
rect 15 -1375 73 -1363
rect 15 -1551 27 -1375
rect 61 -1551 73 -1375
rect 15 -1563 73 -1551
rect -73 -1793 -15 -1781
rect -73 -1969 -61 -1793
rect -27 -1969 -15 -1793
rect -73 -1981 -15 -1969
rect 15 -1793 73 -1781
rect 15 -1969 27 -1793
rect 61 -1969 73 -1793
rect 15 -1981 73 -1969
<< ndiffc >>
rect -61 1793 -27 1969
rect 27 1793 61 1969
rect -61 1375 -27 1551
rect 27 1375 61 1551
rect -61 957 -27 1133
rect 27 957 61 1133
rect -61 539 -27 715
rect 27 539 61 715
rect -61 121 -27 297
rect 27 121 61 297
rect -61 -297 -27 -121
rect 27 -297 61 -121
rect -61 -715 -27 -539
rect 27 -715 61 -539
rect -61 -1133 -27 -957
rect 27 -1133 61 -957
rect -61 -1551 -27 -1375
rect 27 -1551 61 -1375
rect -61 -1969 -27 -1793
rect 27 -1969 61 -1793
<< psubdiff >>
rect -175 2121 -79 2155
rect 79 2121 175 2155
rect -175 2059 -141 2121
rect 141 2059 175 2121
rect -175 -2121 -141 -2059
rect 141 -2121 175 -2059
rect -175 -2155 -79 -2121
rect 79 -2155 175 -2121
<< psubdiffcont >>
rect -79 2121 79 2155
rect -175 -2059 -141 2059
rect 141 -2059 175 2059
rect -79 -2155 79 -2121
<< poly >>
rect -33 2053 33 2069
rect -33 2019 -17 2053
rect 17 2019 33 2053
rect -33 2003 33 2019
rect -15 1981 15 2003
rect -15 1759 15 1781
rect -33 1743 33 1759
rect -33 1709 -17 1743
rect 17 1709 33 1743
rect -33 1693 33 1709
rect -33 1635 33 1651
rect -33 1601 -17 1635
rect 17 1601 33 1635
rect -33 1585 33 1601
rect -15 1563 15 1585
rect -15 1341 15 1363
rect -33 1325 33 1341
rect -33 1291 -17 1325
rect 17 1291 33 1325
rect -33 1275 33 1291
rect -33 1217 33 1233
rect -33 1183 -17 1217
rect 17 1183 33 1217
rect -33 1167 33 1183
rect -15 1145 15 1167
rect -15 923 15 945
rect -33 907 33 923
rect -33 873 -17 907
rect 17 873 33 907
rect -33 857 33 873
rect -33 799 33 815
rect -33 765 -17 799
rect 17 765 33 799
rect -33 749 33 765
rect -15 727 15 749
rect -15 505 15 527
rect -33 489 33 505
rect -33 455 -17 489
rect 17 455 33 489
rect -33 439 33 455
rect -33 381 33 397
rect -33 347 -17 381
rect 17 347 33 381
rect -33 331 33 347
rect -15 309 15 331
rect -15 87 15 109
rect -33 71 33 87
rect -33 37 -17 71
rect 17 37 33 71
rect -33 21 33 37
rect -33 -37 33 -21
rect -33 -71 -17 -37
rect 17 -71 33 -37
rect -33 -87 33 -71
rect -15 -109 15 -87
rect -15 -331 15 -309
rect -33 -347 33 -331
rect -33 -381 -17 -347
rect 17 -381 33 -347
rect -33 -397 33 -381
rect -33 -455 33 -439
rect -33 -489 -17 -455
rect 17 -489 33 -455
rect -33 -505 33 -489
rect -15 -527 15 -505
rect -15 -749 15 -727
rect -33 -765 33 -749
rect -33 -799 -17 -765
rect 17 -799 33 -765
rect -33 -815 33 -799
rect -33 -873 33 -857
rect -33 -907 -17 -873
rect 17 -907 33 -873
rect -33 -923 33 -907
rect -15 -945 15 -923
rect -15 -1167 15 -1145
rect -33 -1183 33 -1167
rect -33 -1217 -17 -1183
rect 17 -1217 33 -1183
rect -33 -1233 33 -1217
rect -33 -1291 33 -1275
rect -33 -1325 -17 -1291
rect 17 -1325 33 -1291
rect -33 -1341 33 -1325
rect -15 -1363 15 -1341
rect -15 -1585 15 -1563
rect -33 -1601 33 -1585
rect -33 -1635 -17 -1601
rect 17 -1635 33 -1601
rect -33 -1651 33 -1635
rect -33 -1709 33 -1693
rect -33 -1743 -17 -1709
rect 17 -1743 33 -1709
rect -33 -1759 33 -1743
rect -15 -1781 15 -1759
rect -15 -2003 15 -1981
rect -33 -2019 33 -2003
rect -33 -2053 -17 -2019
rect 17 -2053 33 -2019
rect -33 -2069 33 -2053
<< polycont >>
rect -17 2019 17 2053
rect -17 1709 17 1743
rect -17 1601 17 1635
rect -17 1291 17 1325
rect -17 1183 17 1217
rect -17 873 17 907
rect -17 765 17 799
rect -17 455 17 489
rect -17 347 17 381
rect -17 37 17 71
rect -17 -71 17 -37
rect -17 -381 17 -347
rect -17 -489 17 -455
rect -17 -799 17 -765
rect -17 -907 17 -873
rect -17 -1217 17 -1183
rect -17 -1325 17 -1291
rect -17 -1635 17 -1601
rect -17 -1743 17 -1709
rect -17 -2053 17 -2019
<< locali >>
rect -175 2121 -79 2155
rect 79 2121 175 2155
rect -175 2059 -141 2121
rect 141 2059 175 2121
rect -33 2019 -17 2053
rect 17 2019 33 2053
rect -61 1969 -27 1985
rect -61 1777 -27 1793
rect 27 1969 61 1985
rect 27 1777 61 1793
rect -33 1709 -17 1743
rect 17 1709 33 1743
rect -33 1601 -17 1635
rect 17 1601 33 1635
rect -61 1551 -27 1567
rect -61 1359 -27 1375
rect 27 1551 61 1567
rect 27 1359 61 1375
rect -33 1291 -17 1325
rect 17 1291 33 1325
rect -33 1183 -17 1217
rect 17 1183 33 1217
rect -61 1133 -27 1149
rect -61 941 -27 957
rect 27 1133 61 1149
rect 27 941 61 957
rect -33 873 -17 907
rect 17 873 33 907
rect -33 765 -17 799
rect 17 765 33 799
rect -61 715 -27 731
rect -61 523 -27 539
rect 27 715 61 731
rect 27 523 61 539
rect -33 455 -17 489
rect 17 455 33 489
rect -33 347 -17 381
rect 17 347 33 381
rect -61 297 -27 313
rect -61 105 -27 121
rect 27 297 61 313
rect 27 105 61 121
rect -33 37 -17 71
rect 17 37 33 71
rect -33 -71 -17 -37
rect 17 -71 33 -37
rect -61 -121 -27 -105
rect -61 -313 -27 -297
rect 27 -121 61 -105
rect 27 -313 61 -297
rect -33 -381 -17 -347
rect 17 -381 33 -347
rect -33 -489 -17 -455
rect 17 -489 33 -455
rect -61 -539 -27 -523
rect -61 -731 -27 -715
rect 27 -539 61 -523
rect 27 -731 61 -715
rect -33 -799 -17 -765
rect 17 -799 33 -765
rect -33 -907 -17 -873
rect 17 -907 33 -873
rect -61 -957 -27 -941
rect -61 -1149 -27 -1133
rect 27 -957 61 -941
rect 27 -1149 61 -1133
rect -33 -1217 -17 -1183
rect 17 -1217 33 -1183
rect -33 -1325 -17 -1291
rect 17 -1325 33 -1291
rect -61 -1375 -27 -1359
rect -61 -1567 -27 -1551
rect 27 -1375 61 -1359
rect 27 -1567 61 -1551
rect -33 -1635 -17 -1601
rect 17 -1635 33 -1601
rect -33 -1743 -17 -1709
rect 17 -1743 33 -1709
rect -61 -1793 -27 -1777
rect -61 -1985 -27 -1969
rect 27 -1793 61 -1777
rect 27 -1985 61 -1969
rect -33 -2053 -17 -2019
rect 17 -2053 33 -2019
rect -175 -2121 -141 -2059
rect 141 -2121 175 -2059
rect -175 -2155 -79 -2121
rect 79 -2155 175 -2121
<< viali >>
rect -17 2019 17 2053
rect -61 1793 -27 1969
rect 27 1793 61 1969
rect -17 1709 17 1743
rect -17 1601 17 1635
rect -61 1375 -27 1551
rect 27 1375 61 1551
rect -17 1291 17 1325
rect -17 1183 17 1217
rect -61 957 -27 1133
rect 27 957 61 1133
rect -17 873 17 907
rect -17 765 17 799
rect -61 539 -27 715
rect 27 539 61 715
rect -17 455 17 489
rect -17 347 17 381
rect -61 121 -27 297
rect 27 121 61 297
rect -17 37 17 71
rect -17 -71 17 -37
rect -61 -297 -27 -121
rect 27 -297 61 -121
rect -17 -381 17 -347
rect -17 -489 17 -455
rect -61 -715 -27 -539
rect 27 -715 61 -539
rect -17 -799 17 -765
rect -17 -907 17 -873
rect -61 -1133 -27 -957
rect 27 -1133 61 -957
rect -17 -1217 17 -1183
rect -17 -1325 17 -1291
rect -61 -1551 -27 -1375
rect 27 -1551 61 -1375
rect -17 -1635 17 -1601
rect -17 -1743 17 -1709
rect -61 -1969 -27 -1793
rect 27 -1969 61 -1793
rect -17 -2053 17 -2019
<< metal1 >>
rect -29 2053 29 2059
rect -29 2019 -17 2053
rect 17 2019 29 2053
rect -29 2013 29 2019
rect -67 1969 -21 1981
rect -67 1793 -61 1969
rect -27 1793 -21 1969
rect -67 1781 -21 1793
rect 21 1969 67 1981
rect 21 1793 27 1969
rect 61 1793 67 1969
rect 21 1781 67 1793
rect -29 1743 29 1749
rect -29 1709 -17 1743
rect 17 1709 29 1743
rect -29 1703 29 1709
rect -29 1635 29 1641
rect -29 1601 -17 1635
rect 17 1601 29 1635
rect -29 1595 29 1601
rect -67 1551 -21 1563
rect -67 1375 -61 1551
rect -27 1375 -21 1551
rect -67 1363 -21 1375
rect 21 1551 67 1563
rect 21 1375 27 1551
rect 61 1375 67 1551
rect 21 1363 67 1375
rect -29 1325 29 1331
rect -29 1291 -17 1325
rect 17 1291 29 1325
rect -29 1285 29 1291
rect -29 1217 29 1223
rect -29 1183 -17 1217
rect 17 1183 29 1217
rect -29 1177 29 1183
rect -67 1133 -21 1145
rect -67 957 -61 1133
rect -27 957 -21 1133
rect -67 945 -21 957
rect 21 1133 67 1145
rect 21 957 27 1133
rect 61 957 67 1133
rect 21 945 67 957
rect -29 907 29 913
rect -29 873 -17 907
rect 17 873 29 907
rect -29 867 29 873
rect -29 799 29 805
rect -29 765 -17 799
rect 17 765 29 799
rect -29 759 29 765
rect -67 715 -21 727
rect -67 539 -61 715
rect -27 539 -21 715
rect -67 527 -21 539
rect 21 715 67 727
rect 21 539 27 715
rect 61 539 67 715
rect 21 527 67 539
rect -29 489 29 495
rect -29 455 -17 489
rect 17 455 29 489
rect -29 449 29 455
rect -29 381 29 387
rect -29 347 -17 381
rect 17 347 29 381
rect -29 341 29 347
rect -67 297 -21 309
rect -67 121 -61 297
rect -27 121 -21 297
rect -67 109 -21 121
rect 21 297 67 309
rect 21 121 27 297
rect 61 121 67 297
rect 21 109 67 121
rect -29 71 29 77
rect -29 37 -17 71
rect 17 37 29 71
rect -29 31 29 37
rect -29 -37 29 -31
rect -29 -71 -17 -37
rect 17 -71 29 -37
rect -29 -77 29 -71
rect -67 -121 -21 -109
rect -67 -297 -61 -121
rect -27 -297 -21 -121
rect -67 -309 -21 -297
rect 21 -121 67 -109
rect 21 -297 27 -121
rect 61 -297 67 -121
rect 21 -309 67 -297
rect -29 -347 29 -341
rect -29 -381 -17 -347
rect 17 -381 29 -347
rect -29 -387 29 -381
rect -29 -455 29 -449
rect -29 -489 -17 -455
rect 17 -489 29 -455
rect -29 -495 29 -489
rect -67 -539 -21 -527
rect -67 -715 -61 -539
rect -27 -715 -21 -539
rect -67 -727 -21 -715
rect 21 -539 67 -527
rect 21 -715 27 -539
rect 61 -715 67 -539
rect 21 -727 67 -715
rect -29 -765 29 -759
rect -29 -799 -17 -765
rect 17 -799 29 -765
rect -29 -805 29 -799
rect -29 -873 29 -867
rect -29 -907 -17 -873
rect 17 -907 29 -873
rect -29 -913 29 -907
rect -67 -957 -21 -945
rect -67 -1133 -61 -957
rect -27 -1133 -21 -957
rect -67 -1145 -21 -1133
rect 21 -957 67 -945
rect 21 -1133 27 -957
rect 61 -1133 67 -957
rect 21 -1145 67 -1133
rect -29 -1183 29 -1177
rect -29 -1217 -17 -1183
rect 17 -1217 29 -1183
rect -29 -1223 29 -1217
rect -29 -1291 29 -1285
rect -29 -1325 -17 -1291
rect 17 -1325 29 -1291
rect -29 -1331 29 -1325
rect -67 -1375 -21 -1363
rect -67 -1551 -61 -1375
rect -27 -1551 -21 -1375
rect -67 -1563 -21 -1551
rect 21 -1375 67 -1363
rect 21 -1551 27 -1375
rect 61 -1551 67 -1375
rect 21 -1563 67 -1551
rect -29 -1601 29 -1595
rect -29 -1635 -17 -1601
rect 17 -1635 29 -1601
rect -29 -1641 29 -1635
rect -29 -1709 29 -1703
rect -29 -1743 -17 -1709
rect 17 -1743 29 -1709
rect -29 -1749 29 -1743
rect -67 -1793 -21 -1781
rect -67 -1969 -61 -1793
rect -27 -1969 -21 -1793
rect -67 -1981 -21 -1969
rect 21 -1793 67 -1781
rect 21 -1969 27 -1793
rect 61 -1969 67 -1793
rect 21 -1981 67 -1969
rect -29 -2019 29 -2013
rect -29 -2053 -17 -2019
rect 17 -2053 29 -2019
rect -29 -2059 29 -2053
<< properties >>
string FIXED_BBOX -158 -2138 158 2138
string gencell sky130_fd_pr__nfet_01v8_lvt
string library sky130
string parameters w 1 l 0.150 m 10 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
