magic
tech sky130A
magscale 1 2
timestamp 1672277640
<< locali >>
rect 180 360 240 540
rect 1100 360 1160 540
rect 2020 360 2080 540
rect 2920 360 2980 540
rect 3840 360 3900 540
rect 4760 360 4820 540
rect 5220 360 5280 540
<< metal1 >>
rect 1050 7820 1060 7920
rect 1160 7820 1170 7920
rect 1970 7820 1980 7920
rect 2080 7820 2090 7920
rect 2890 7820 2900 7920
rect 3000 7820 3010 7920
rect 3810 7820 3820 7920
rect 3920 7820 3930 7920
rect 4730 7820 4740 7920
rect 4840 7820 4850 7920
rect 1510 6800 1520 6900
rect 1620 6800 1630 6900
rect 4270 6800 4280 6900
rect 4380 6800 4390 6900
rect 2430 5600 2440 5700
rect 2540 5600 2550 5700
rect 3350 5600 3360 5700
rect 3460 5600 3470 5700
rect 1520 4630 4520 4780
rect 2430 3700 2440 3800
rect 2540 3700 2550 3800
rect 3350 3700 3360 3800
rect 3460 3700 3470 3800
rect 1510 2600 1520 2700
rect 1620 2600 1630 2700
rect 4270 2600 4280 2700
rect 4390 2600 4400 2700
rect 1070 1480 1080 1580
rect 1180 1480 1190 1580
rect 1970 1480 1980 1580
rect 2080 1480 2090 1580
rect 2890 1480 2900 1580
rect 3000 1480 3010 1580
rect 3810 1480 3820 1580
rect 3920 1480 3930 1580
rect 4730 1480 4740 1580
rect 4840 1480 4850 1580
rect 180 160 280 900
rect 1080 870 4380 900
rect 1070 700 1080 780
rect 1160 700 1170 780
rect 1990 700 2000 780
rect 2080 700 2090 780
rect 2910 700 2920 780
rect 3000 700 3010 780
rect 3810 700 3820 780
rect 3900 700 3910 780
rect 4730 700 4740 780
rect 4820 700 4830 780
rect 640 580 700 680
rect 1560 580 1620 680
rect 2480 580 2540 680
rect 3380 580 3440 680
rect 4300 580 4360 680
rect 640 480 4360 580
rect 640 380 700 480
rect 1560 380 1620 480
rect 2480 380 2540 480
rect 3380 380 3440 480
rect 4300 380 4360 480
rect 1080 160 4380 190
rect 5160 160 5280 920
<< via1 >>
rect 1060 7820 1160 7920
rect 1980 7820 2080 7920
rect 2900 7820 3000 7920
rect 3820 7820 3920 7920
rect 4740 7820 4840 7920
rect 1520 6800 1620 6900
rect 4280 6800 4380 6900
rect 2440 5600 2540 5700
rect 3360 5600 3460 5700
rect 2440 3700 2540 3800
rect 3360 3700 3460 3800
rect 1520 2600 1620 2700
rect 4280 2600 4390 2700
rect 1080 1480 1180 1580
rect 1980 1480 2080 1580
rect 2900 1480 3000 1580
rect 3820 1480 3920 1580
rect 4740 1480 4840 1580
rect 1080 700 1160 780
rect 2000 700 2080 780
rect 2920 700 3000 780
rect 3820 700 3900 780
rect 4740 700 4820 780
<< metal2 >>
rect 1060 7920 4840 7940
rect 1160 7820 1980 7920
rect 2080 7820 2900 7920
rect 3000 7820 3820 7920
rect 3920 7820 4740 7920
rect 1060 7800 4840 7820
rect 1500 6900 4400 6920
rect 1500 6800 1520 6900
rect 1620 6800 4280 6900
rect 4380 6800 4400 6900
rect 1500 6780 4400 6800
rect 1500 5700 3460 5720
rect 1500 5600 2440 5700
rect 2540 5600 3360 5700
rect 1500 5580 3460 5600
rect 1500 2720 1640 5580
rect 4260 3820 4400 6780
rect 2440 3800 4400 3820
rect 2540 3700 3360 3800
rect 3460 3700 4400 3800
rect 2440 3680 4400 3700
rect 1500 2700 4400 2720
rect 1500 2600 1520 2700
rect 1620 2600 2800 2700
rect 1500 2580 2800 2600
rect 3100 2600 4280 2700
rect 4390 2600 4400 2700
rect 3100 2580 4400 2600
rect 2800 2490 3100 2500
rect 1080 1580 4840 1600
rect 1180 1480 1980 1580
rect 2080 1480 2900 1580
rect 3000 1480 3820 1580
rect 3920 1480 4740 1580
rect 1080 1460 4840 1480
rect 2800 800 3100 810
rect 1080 780 1160 790
rect 2000 780 2080 790
rect 3820 780 3900 790
rect 4740 780 4820 790
rect 1060 700 1080 780
rect 1160 700 2000 780
rect 2080 700 2800 780
rect 3100 700 3820 780
rect 3900 700 4740 780
rect 4820 700 4840 780
rect 1080 690 1160 700
rect 2000 690 2080 700
rect 3820 690 3900 700
rect 4740 690 4820 700
rect 2800 590 3100 600
<< via2 >>
rect 2800 2500 3100 2700
rect 2800 780 3100 800
rect 2800 700 2920 780
rect 2920 700 3000 780
rect 3000 700 3100 780
rect 2800 600 3100 700
<< metal3 >>
rect 2800 2705 3100 2800
rect 2790 2700 3110 2705
rect 2790 2500 2800 2700
rect 3100 2500 3110 2700
rect 2790 2495 3110 2500
rect 2800 805 3100 2495
rect 2790 800 3110 805
rect 2790 600 2800 800
rect 3100 600 3110 800
rect 2790 595 3110 600
use sky130_fd_pr__nfet_01v8_lvt_J9QE6F  sky130_fd_pr__nfet_01v8_lvt_J9QE6F_1
timestamp 1672262880
transform 1 0 2726 0 1 299
box -2686 -279 2686 279
use sky130_fd_pr__nfet_01v8_lvt_M93XMJ  sky130_fd_pr__nfet_01v8_lvt_M93XMJ_0
timestamp 1672262880
transform 1 0 2726 0 1 759
box -2686 -279 2686 279
use sky130_fd_pr__pfet_01v8_lvt_QH9SH3  sky130_fd_pr__pfet_01v8_lvt_QH9SH3_0
timestamp 1672264357
transform 1 0 2723 0 1 4704
box -2686 -3537 2686 3537
<< labels >>
flabel space 1080 -180 1180 -20 0 FreeSans 800 0 0 0 S
flabel space 1980 -160 2080 0 0 FreeSans 800 0 0 0 S
flabel space 2900 -140 3000 20 0 FreeSans 800 0 0 0 S
flabel space 3820 -140 3920 20 0 FreeSans 800 0 0 0 S
flabel space 4740 -160 4840 0 0 FreeSans 800 0 0 0 S
flabel space 1520 -180 1620 -20 0 FreeSans 800 0 0 0 D
flabel space 2440 -180 2540 -20 0 FreeSans 800 0 0 0 D
flabel space 3360 -140 3460 20 0 FreeSans 800 0 0 0 D
flabel space 4280 -120 4380 40 0 FreeSans 800 0 0 0 D
flabel space 620 -200 720 -40 0 FreeSans 800 0 0 0 D
flabel space 1280 1030 1380 1180 0 FreeSans 800 0 0 0 A
flabel space 1760 1030 1860 1180 0 FreeSans 800 0 0 0 A
flabel space 4030 1060 4130 1210 0 FreeSans 800 0 0 0 A
flabel space 4520 1050 4620 1200 0 FreeSans 800 0 0 0 A
flabel space 2220 1030 2320 1180 0 FreeSans 800 0 0 0 B
flabel space 2690 1020 2790 1170 0 FreeSans 800 0 0 0 B
flabel space 3130 1010 3230 1160 0 FreeSans 800 0 0 0 B
flabel space 3580 1040 3680 1190 0 FreeSans 800 0 0 0 B
flabel space 1290 8290 1390 8440 0 FreeSans 800 0 0 0 B
flabel space 1730 8290 1830 8440 0 FreeSans 800 0 0 0 B
flabel space 2210 8290 2310 8440 0 FreeSans 800 0 0 0 A
flabel space 2660 8300 2760 8450 0 FreeSans 800 0 0 0 A
flabel space 3110 8280 3210 8430 0 FreeSans 800 0 0 0 A
flabel space 3590 8290 3690 8440 0 FreeSans 800 0 0 0 A
flabel space 4060 8280 4160 8430 0 FreeSans 800 0 0 0 B
flabel space 4530 8280 4630 8430 0 FreeSans 800 0 0 0 B
<< end >>
