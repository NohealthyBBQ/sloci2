magic
tech sky130A
magscale 1 2
timestamp 1672262786
<< pwell >>
rect -2228 -279 2228 279
<< nmoslvt >>
rect -2032 -69 -1632 131
rect -1574 -69 -1174 131
rect -1116 -69 -716 131
rect -658 -69 -258 131
rect -200 -69 200 131
rect 258 -69 658 131
rect 716 -69 1116 131
rect 1174 -69 1574 131
rect 1632 -69 2032 131
<< ndiff >>
rect -2090 119 -2032 131
rect -2090 -57 -2078 119
rect -2044 -57 -2032 119
rect -2090 -69 -2032 -57
rect -1632 119 -1574 131
rect -1632 -57 -1620 119
rect -1586 -57 -1574 119
rect -1632 -69 -1574 -57
rect -1174 119 -1116 131
rect -1174 -57 -1162 119
rect -1128 -57 -1116 119
rect -1174 -69 -1116 -57
rect -716 119 -658 131
rect -716 -57 -704 119
rect -670 -57 -658 119
rect -716 -69 -658 -57
rect -258 119 -200 131
rect -258 -57 -246 119
rect -212 -57 -200 119
rect -258 -69 -200 -57
rect 200 119 258 131
rect 200 -57 212 119
rect 246 -57 258 119
rect 200 -69 258 -57
rect 658 119 716 131
rect 658 -57 670 119
rect 704 -57 716 119
rect 658 -69 716 -57
rect 1116 119 1174 131
rect 1116 -57 1128 119
rect 1162 -57 1174 119
rect 1116 -69 1174 -57
rect 1574 119 1632 131
rect 1574 -57 1586 119
rect 1620 -57 1632 119
rect 1574 -69 1632 -57
rect 2032 119 2090 131
rect 2032 -57 2044 119
rect 2078 -57 2090 119
rect 2032 -69 2090 -57
<< ndiffc >>
rect -2078 -57 -2044 119
rect -1620 -57 -1586 119
rect -1162 -57 -1128 119
rect -704 -57 -670 119
rect -246 -57 -212 119
rect 212 -57 246 119
rect 670 -57 704 119
rect 1128 -57 1162 119
rect 1586 -57 1620 119
rect 2044 -57 2078 119
<< psubdiff >>
rect -2192 209 2192 243
rect -2192 -209 -2158 209
rect 2158 -209 2192 209
rect -2192 -243 -2096 -209
rect 2096 -243 2192 -209
<< psubdiffcont >>
rect -2096 -243 2096 -209
<< poly >>
rect -2032 131 -1632 157
rect -1574 131 -1174 157
rect -1116 131 -716 157
rect -658 131 -258 157
rect -200 131 200 157
rect 258 131 658 157
rect 716 131 1116 157
rect 1174 131 1574 157
rect 1632 131 2032 157
rect -2032 -107 -1632 -69
rect -2032 -141 -2016 -107
rect -1648 -141 -1632 -107
rect -2032 -157 -1632 -141
rect -1574 -107 -1174 -69
rect -1574 -141 -1558 -107
rect -1190 -141 -1174 -107
rect -1574 -157 -1174 -141
rect -1116 -107 -716 -69
rect -1116 -141 -1100 -107
rect -732 -141 -716 -107
rect -1116 -157 -716 -141
rect -658 -107 -258 -69
rect -658 -141 -642 -107
rect -274 -141 -258 -107
rect -658 -157 -258 -141
rect -200 -107 200 -69
rect -200 -141 -184 -107
rect 184 -141 200 -107
rect -200 -157 200 -141
rect 258 -107 658 -69
rect 258 -141 274 -107
rect 642 -141 658 -107
rect 258 -157 658 -141
rect 716 -107 1116 -69
rect 716 -141 732 -107
rect 1100 -141 1116 -107
rect 716 -157 1116 -141
rect 1174 -107 1574 -69
rect 1174 -141 1190 -107
rect 1558 -141 1574 -107
rect 1174 -157 1574 -141
rect 1632 -107 2032 -69
rect 1632 -141 1648 -107
rect 2016 -141 2032 -107
rect 1632 -157 2032 -141
<< polycont >>
rect -2016 -141 -1648 -107
rect -1558 -141 -1190 -107
rect -1100 -141 -732 -107
rect -642 -141 -274 -107
rect -184 -141 184 -107
rect 274 -141 642 -107
rect 732 -141 1100 -107
rect 1190 -141 1558 -107
rect 1648 -141 2016 -107
<< locali >>
rect -2192 209 2192 243
rect -2192 -209 -2158 209
rect -2078 119 -2044 135
rect -2078 -73 -2044 -57
rect -1620 119 -1586 135
rect -1620 -73 -1586 -57
rect -1162 119 -1128 135
rect -1162 -73 -1128 -57
rect -704 119 -670 135
rect -704 -73 -670 -57
rect -246 119 -212 135
rect -246 -73 -212 -57
rect 212 119 246 135
rect 212 -73 246 -57
rect 670 119 704 135
rect 670 -73 704 -57
rect 1128 119 1162 135
rect 1128 -73 1162 -57
rect 1586 119 1620 135
rect 1586 -73 1620 -57
rect 2044 119 2078 135
rect 2044 -73 2078 -57
rect -2032 -141 -2016 -107
rect -1648 -141 -1632 -107
rect -1574 -141 -1558 -107
rect -1190 -141 -1174 -107
rect -1116 -141 -1100 -107
rect -732 -141 -716 -107
rect -658 -141 -642 -107
rect -274 -141 -258 -107
rect -200 -141 -184 -107
rect 184 -141 200 -107
rect 258 -141 274 -107
rect 642 -141 658 -107
rect 716 -141 732 -107
rect 1100 -141 1116 -107
rect 1174 -141 1190 -107
rect 1558 -141 1574 -107
rect 1632 -141 1648 -107
rect 2016 -141 2032 -107
rect 2158 -209 2192 209
rect -2192 -243 -2096 -209
rect 2096 -243 2192 -209
<< viali >>
rect -2078 -57 -2044 119
rect -1620 -57 -1586 119
rect -1162 -57 -1128 119
rect -704 -57 -670 119
rect -246 -57 -212 119
rect 212 -57 246 119
rect 670 -57 704 119
rect 1128 -57 1162 119
rect 1586 -57 1620 119
rect 2044 -57 2078 119
rect -2016 -141 -1648 -107
rect -1558 -141 -1190 -107
rect -1100 -141 -732 -107
rect -642 -141 -274 -107
rect -184 -141 184 -107
rect 274 -141 642 -107
rect 732 -141 1100 -107
rect 1190 -141 1558 -107
rect 1648 -141 2016 -107
<< metal1 >>
rect -2084 119 -2038 131
rect -2084 -57 -2078 119
rect -2044 -57 -2038 119
rect -2084 -69 -2038 -57
rect -1626 119 -1580 131
rect -1626 -57 -1620 119
rect -1586 -57 -1580 119
rect -1626 -69 -1580 -57
rect -1168 119 -1122 131
rect -1168 -57 -1162 119
rect -1128 -57 -1122 119
rect -1168 -69 -1122 -57
rect -710 119 -664 131
rect -710 -57 -704 119
rect -670 -57 -664 119
rect -710 -69 -664 -57
rect -252 119 -206 131
rect -252 -57 -246 119
rect -212 -57 -206 119
rect -252 -69 -206 -57
rect 206 119 252 131
rect 206 -57 212 119
rect 246 -57 252 119
rect 206 -69 252 -57
rect 664 119 710 131
rect 664 -57 670 119
rect 704 -57 710 119
rect 664 -69 710 -57
rect 1122 119 1168 131
rect 1122 -57 1128 119
rect 1162 -57 1168 119
rect 1122 -69 1168 -57
rect 1580 119 1626 131
rect 1580 -57 1586 119
rect 1620 -57 1626 119
rect 1580 -69 1626 -57
rect 2038 119 2084 131
rect 2038 -57 2044 119
rect 2078 -57 2084 119
rect 2038 -69 2084 -57
rect -2028 -107 -1636 -101
rect -2028 -141 -2016 -107
rect -1648 -141 -1636 -107
rect -2028 -147 -1636 -141
rect -1570 -107 -1178 -101
rect -1570 -141 -1558 -107
rect -1190 -141 -1178 -107
rect -1570 -147 -1178 -141
rect -1112 -107 -720 -101
rect -1112 -141 -1100 -107
rect -732 -141 -720 -107
rect -1112 -147 -720 -141
rect -654 -107 -262 -101
rect -654 -141 -642 -107
rect -274 -141 -262 -107
rect -654 -147 -262 -141
rect -196 -107 196 -101
rect -196 -141 -184 -107
rect 184 -141 196 -107
rect -196 -147 196 -141
rect 262 -107 654 -101
rect 262 -141 274 -107
rect 642 -141 654 -107
rect 262 -147 654 -141
rect 720 -107 1112 -101
rect 720 -141 732 -107
rect 1100 -141 1112 -107
rect 720 -147 1112 -141
rect 1178 -107 1570 -101
rect 1178 -141 1190 -107
rect 1558 -141 1570 -107
rect 1178 -147 1570 -141
rect 1636 -107 2028 -101
rect 1636 -141 1648 -107
rect 2016 -141 2028 -107
rect 1636 -147 2028 -141
<< properties >>
string FIXED_BBOX -2175 -226 2175 226
string gencell sky130_fd_pr__nfet_01v8_lvt
string library sky130
string parameters w 1 l 2 m 1 nf 9 diffcov 100 polycov 100 guard 1 glc 0 grc 0 gtc 0 gbc 1 tbcov 100 rlcov 100 topc 0 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
