magic
tech sky130A
magscale 1 2
timestamp 1662478139
<< pwell >>
rect -396 -2191 396 2191
<< nmoslvt >>
rect -200 1781 200 1981
rect -200 1363 200 1563
rect -200 945 200 1145
rect -200 527 200 727
rect -200 109 200 309
rect -200 -309 200 -109
rect -200 -727 200 -527
rect -200 -1145 200 -945
rect -200 -1563 200 -1363
rect -200 -1981 200 -1781
<< ndiff >>
rect -258 1969 -200 1981
rect -258 1793 -246 1969
rect -212 1793 -200 1969
rect -258 1781 -200 1793
rect 200 1969 258 1981
rect 200 1793 212 1969
rect 246 1793 258 1969
rect 200 1781 258 1793
rect -258 1551 -200 1563
rect -258 1375 -246 1551
rect -212 1375 -200 1551
rect -258 1363 -200 1375
rect 200 1551 258 1563
rect 200 1375 212 1551
rect 246 1375 258 1551
rect 200 1363 258 1375
rect -258 1133 -200 1145
rect -258 957 -246 1133
rect -212 957 -200 1133
rect -258 945 -200 957
rect 200 1133 258 1145
rect 200 957 212 1133
rect 246 957 258 1133
rect 200 945 258 957
rect -258 715 -200 727
rect -258 539 -246 715
rect -212 539 -200 715
rect -258 527 -200 539
rect 200 715 258 727
rect 200 539 212 715
rect 246 539 258 715
rect 200 527 258 539
rect -258 297 -200 309
rect -258 121 -246 297
rect -212 121 -200 297
rect -258 109 -200 121
rect 200 297 258 309
rect 200 121 212 297
rect 246 121 258 297
rect 200 109 258 121
rect -258 -121 -200 -109
rect -258 -297 -246 -121
rect -212 -297 -200 -121
rect -258 -309 -200 -297
rect 200 -121 258 -109
rect 200 -297 212 -121
rect 246 -297 258 -121
rect 200 -309 258 -297
rect -258 -539 -200 -527
rect -258 -715 -246 -539
rect -212 -715 -200 -539
rect -258 -727 -200 -715
rect 200 -539 258 -527
rect 200 -715 212 -539
rect 246 -715 258 -539
rect 200 -727 258 -715
rect -258 -957 -200 -945
rect -258 -1133 -246 -957
rect -212 -1133 -200 -957
rect -258 -1145 -200 -1133
rect 200 -957 258 -945
rect 200 -1133 212 -957
rect 246 -1133 258 -957
rect 200 -1145 258 -1133
rect -258 -1375 -200 -1363
rect -258 -1551 -246 -1375
rect -212 -1551 -200 -1375
rect -258 -1563 -200 -1551
rect 200 -1375 258 -1363
rect 200 -1551 212 -1375
rect 246 -1551 258 -1375
rect 200 -1563 258 -1551
rect -258 -1793 -200 -1781
rect -258 -1969 -246 -1793
rect -212 -1969 -200 -1793
rect -258 -1981 -200 -1969
rect 200 -1793 258 -1781
rect 200 -1969 212 -1793
rect 246 -1969 258 -1793
rect 200 -1981 258 -1969
<< ndiffc >>
rect -246 1793 -212 1969
rect 212 1793 246 1969
rect -246 1375 -212 1551
rect 212 1375 246 1551
rect -246 957 -212 1133
rect 212 957 246 1133
rect -246 539 -212 715
rect 212 539 246 715
rect -246 121 -212 297
rect 212 121 246 297
rect -246 -297 -212 -121
rect 212 -297 246 -121
rect -246 -715 -212 -539
rect 212 -715 246 -539
rect -246 -1133 -212 -957
rect 212 -1133 246 -957
rect -246 -1551 -212 -1375
rect 212 -1551 246 -1375
rect -246 -1969 -212 -1793
rect 212 -1969 246 -1793
<< psubdiff >>
rect -360 2121 -264 2155
rect 264 2121 360 2155
rect -360 2059 -326 2121
rect 326 2059 360 2121
rect -360 -2121 -326 -2059
rect 326 -2121 360 -2059
rect -360 -2155 -264 -2121
rect 264 -2155 360 -2121
<< psubdiffcont >>
rect -264 2121 264 2155
rect -360 -2059 -326 2059
rect 326 -2059 360 2059
rect -264 -2155 264 -2121
<< poly >>
rect -200 2053 200 2069
rect -200 2019 -184 2053
rect 184 2019 200 2053
rect -200 1981 200 2019
rect -200 1743 200 1781
rect -200 1709 -184 1743
rect 184 1709 200 1743
rect -200 1693 200 1709
rect -200 1635 200 1651
rect -200 1601 -184 1635
rect 184 1601 200 1635
rect -200 1563 200 1601
rect -200 1325 200 1363
rect -200 1291 -184 1325
rect 184 1291 200 1325
rect -200 1275 200 1291
rect -200 1217 200 1233
rect -200 1183 -184 1217
rect 184 1183 200 1217
rect -200 1145 200 1183
rect -200 907 200 945
rect -200 873 -184 907
rect 184 873 200 907
rect -200 857 200 873
rect -200 799 200 815
rect -200 765 -184 799
rect 184 765 200 799
rect -200 727 200 765
rect -200 489 200 527
rect -200 455 -184 489
rect 184 455 200 489
rect -200 439 200 455
rect -200 381 200 397
rect -200 347 -184 381
rect 184 347 200 381
rect -200 309 200 347
rect -200 71 200 109
rect -200 37 -184 71
rect 184 37 200 71
rect -200 21 200 37
rect -200 -37 200 -21
rect -200 -71 -184 -37
rect 184 -71 200 -37
rect -200 -109 200 -71
rect -200 -347 200 -309
rect -200 -381 -184 -347
rect 184 -381 200 -347
rect -200 -397 200 -381
rect -200 -455 200 -439
rect -200 -489 -184 -455
rect 184 -489 200 -455
rect -200 -527 200 -489
rect -200 -765 200 -727
rect -200 -799 -184 -765
rect 184 -799 200 -765
rect -200 -815 200 -799
rect -200 -873 200 -857
rect -200 -907 -184 -873
rect 184 -907 200 -873
rect -200 -945 200 -907
rect -200 -1183 200 -1145
rect -200 -1217 -184 -1183
rect 184 -1217 200 -1183
rect -200 -1233 200 -1217
rect -200 -1291 200 -1275
rect -200 -1325 -184 -1291
rect 184 -1325 200 -1291
rect -200 -1363 200 -1325
rect -200 -1601 200 -1563
rect -200 -1635 -184 -1601
rect 184 -1635 200 -1601
rect -200 -1651 200 -1635
rect -200 -1709 200 -1693
rect -200 -1743 -184 -1709
rect 184 -1743 200 -1709
rect -200 -1781 200 -1743
rect -200 -2019 200 -1981
rect -200 -2053 -184 -2019
rect 184 -2053 200 -2019
rect -200 -2069 200 -2053
<< polycont >>
rect -184 2019 184 2053
rect -184 1709 184 1743
rect -184 1601 184 1635
rect -184 1291 184 1325
rect -184 1183 184 1217
rect -184 873 184 907
rect -184 765 184 799
rect -184 455 184 489
rect -184 347 184 381
rect -184 37 184 71
rect -184 -71 184 -37
rect -184 -381 184 -347
rect -184 -489 184 -455
rect -184 -799 184 -765
rect -184 -907 184 -873
rect -184 -1217 184 -1183
rect -184 -1325 184 -1291
rect -184 -1635 184 -1601
rect -184 -1743 184 -1709
rect -184 -2053 184 -2019
<< locali >>
rect -360 2121 -264 2155
rect 264 2121 360 2155
rect -360 2059 -326 2121
rect 326 2059 360 2121
rect -200 2019 -184 2053
rect 184 2019 200 2053
rect -246 1969 -212 1985
rect -246 1777 -212 1793
rect 212 1969 246 1985
rect 212 1777 246 1793
rect -200 1709 -184 1743
rect 184 1709 200 1743
rect -200 1601 -184 1635
rect 184 1601 200 1635
rect -246 1551 -212 1567
rect -246 1359 -212 1375
rect 212 1551 246 1567
rect 212 1359 246 1375
rect -200 1291 -184 1325
rect 184 1291 200 1325
rect -200 1183 -184 1217
rect 184 1183 200 1217
rect -246 1133 -212 1149
rect -246 941 -212 957
rect 212 1133 246 1149
rect 212 941 246 957
rect -200 873 -184 907
rect 184 873 200 907
rect -200 765 -184 799
rect 184 765 200 799
rect -246 715 -212 731
rect -246 523 -212 539
rect 212 715 246 731
rect 212 523 246 539
rect -200 455 -184 489
rect 184 455 200 489
rect -200 347 -184 381
rect 184 347 200 381
rect -246 297 -212 313
rect -246 105 -212 121
rect 212 297 246 313
rect 212 105 246 121
rect -200 37 -184 71
rect 184 37 200 71
rect -200 -71 -184 -37
rect 184 -71 200 -37
rect -246 -121 -212 -105
rect -246 -313 -212 -297
rect 212 -121 246 -105
rect 212 -313 246 -297
rect -200 -381 -184 -347
rect 184 -381 200 -347
rect -200 -489 -184 -455
rect 184 -489 200 -455
rect -246 -539 -212 -523
rect -246 -731 -212 -715
rect 212 -539 246 -523
rect 212 -731 246 -715
rect -200 -799 -184 -765
rect 184 -799 200 -765
rect -200 -907 -184 -873
rect 184 -907 200 -873
rect -246 -957 -212 -941
rect -246 -1149 -212 -1133
rect 212 -957 246 -941
rect 212 -1149 246 -1133
rect -200 -1217 -184 -1183
rect 184 -1217 200 -1183
rect -200 -1325 -184 -1291
rect 184 -1325 200 -1291
rect -246 -1375 -212 -1359
rect -246 -1567 -212 -1551
rect 212 -1375 246 -1359
rect 212 -1567 246 -1551
rect -200 -1635 -184 -1601
rect 184 -1635 200 -1601
rect -200 -1743 -184 -1709
rect 184 -1743 200 -1709
rect -246 -1793 -212 -1777
rect -246 -1985 -212 -1969
rect 212 -1793 246 -1777
rect 212 -1985 246 -1969
rect -200 -2053 -184 -2019
rect 184 -2053 200 -2019
rect -360 -2121 -326 -2059
rect 326 -2121 360 -2059
rect -360 -2155 -264 -2121
rect 264 -2155 360 -2121
<< viali >>
rect -184 2019 184 2053
rect -246 1793 -212 1969
rect 212 1793 246 1969
rect -184 1709 184 1743
rect -184 1601 184 1635
rect -246 1375 -212 1551
rect 212 1375 246 1551
rect -184 1291 184 1325
rect -184 1183 184 1217
rect -246 957 -212 1133
rect 212 957 246 1133
rect -184 873 184 907
rect -184 765 184 799
rect -246 539 -212 715
rect 212 539 246 715
rect -184 455 184 489
rect -184 347 184 381
rect -246 121 -212 297
rect 212 121 246 297
rect -184 37 184 71
rect -184 -71 184 -37
rect -246 -297 -212 -121
rect 212 -297 246 -121
rect -184 -381 184 -347
rect -184 -489 184 -455
rect -246 -715 -212 -539
rect 212 -715 246 -539
rect -184 -799 184 -765
rect -184 -907 184 -873
rect -246 -1133 -212 -957
rect 212 -1133 246 -957
rect -184 -1217 184 -1183
rect -184 -1325 184 -1291
rect -246 -1551 -212 -1375
rect 212 -1551 246 -1375
rect -184 -1635 184 -1601
rect -184 -1743 184 -1709
rect -246 -1969 -212 -1793
rect 212 -1969 246 -1793
rect -184 -2053 184 -2019
<< metal1 >>
rect -196 2053 196 2059
rect -196 2019 -184 2053
rect 184 2019 196 2053
rect -196 2013 196 2019
rect -252 1969 -206 1981
rect -252 1793 -246 1969
rect -212 1793 -206 1969
rect -252 1781 -206 1793
rect 206 1969 252 1981
rect 206 1793 212 1969
rect 246 1793 252 1969
rect 206 1781 252 1793
rect -196 1743 196 1749
rect -196 1709 -184 1743
rect 184 1709 196 1743
rect -196 1703 196 1709
rect -196 1635 196 1641
rect -196 1601 -184 1635
rect 184 1601 196 1635
rect -196 1595 196 1601
rect -252 1551 -206 1563
rect -252 1375 -246 1551
rect -212 1375 -206 1551
rect -252 1363 -206 1375
rect 206 1551 252 1563
rect 206 1375 212 1551
rect 246 1375 252 1551
rect 206 1363 252 1375
rect -196 1325 196 1331
rect -196 1291 -184 1325
rect 184 1291 196 1325
rect -196 1285 196 1291
rect -196 1217 196 1223
rect -196 1183 -184 1217
rect 184 1183 196 1217
rect -196 1177 196 1183
rect -252 1133 -206 1145
rect -252 957 -246 1133
rect -212 957 -206 1133
rect -252 945 -206 957
rect 206 1133 252 1145
rect 206 957 212 1133
rect 246 957 252 1133
rect 206 945 252 957
rect -196 907 196 913
rect -196 873 -184 907
rect 184 873 196 907
rect -196 867 196 873
rect -196 799 196 805
rect -196 765 -184 799
rect 184 765 196 799
rect -196 759 196 765
rect -252 715 -206 727
rect -252 539 -246 715
rect -212 539 -206 715
rect -252 527 -206 539
rect 206 715 252 727
rect 206 539 212 715
rect 246 539 252 715
rect 206 527 252 539
rect -196 489 196 495
rect -196 455 -184 489
rect 184 455 196 489
rect -196 449 196 455
rect -196 381 196 387
rect -196 347 -184 381
rect 184 347 196 381
rect -196 341 196 347
rect -252 297 -206 309
rect -252 121 -246 297
rect -212 121 -206 297
rect -252 109 -206 121
rect 206 297 252 309
rect 206 121 212 297
rect 246 121 252 297
rect 206 109 252 121
rect -196 71 196 77
rect -196 37 -184 71
rect 184 37 196 71
rect -196 31 196 37
rect -196 -37 196 -31
rect -196 -71 -184 -37
rect 184 -71 196 -37
rect -196 -77 196 -71
rect -252 -121 -206 -109
rect -252 -297 -246 -121
rect -212 -297 -206 -121
rect -252 -309 -206 -297
rect 206 -121 252 -109
rect 206 -297 212 -121
rect 246 -297 252 -121
rect 206 -309 252 -297
rect -196 -347 196 -341
rect -196 -381 -184 -347
rect 184 -381 196 -347
rect -196 -387 196 -381
rect -196 -455 196 -449
rect -196 -489 -184 -455
rect 184 -489 196 -455
rect -196 -495 196 -489
rect -252 -539 -206 -527
rect -252 -715 -246 -539
rect -212 -715 -206 -539
rect -252 -727 -206 -715
rect 206 -539 252 -527
rect 206 -715 212 -539
rect 246 -715 252 -539
rect 206 -727 252 -715
rect -196 -765 196 -759
rect -196 -799 -184 -765
rect 184 -799 196 -765
rect -196 -805 196 -799
rect -196 -873 196 -867
rect -196 -907 -184 -873
rect 184 -907 196 -873
rect -196 -913 196 -907
rect -252 -957 -206 -945
rect -252 -1133 -246 -957
rect -212 -1133 -206 -957
rect -252 -1145 -206 -1133
rect 206 -957 252 -945
rect 206 -1133 212 -957
rect 246 -1133 252 -957
rect 206 -1145 252 -1133
rect -196 -1183 196 -1177
rect -196 -1217 -184 -1183
rect 184 -1217 196 -1183
rect -196 -1223 196 -1217
rect -196 -1291 196 -1285
rect -196 -1325 -184 -1291
rect 184 -1325 196 -1291
rect -196 -1331 196 -1325
rect -252 -1375 -206 -1363
rect -252 -1551 -246 -1375
rect -212 -1551 -206 -1375
rect -252 -1563 -206 -1551
rect 206 -1375 252 -1363
rect 206 -1551 212 -1375
rect 246 -1551 252 -1375
rect 206 -1563 252 -1551
rect -196 -1601 196 -1595
rect -196 -1635 -184 -1601
rect 184 -1635 196 -1601
rect -196 -1641 196 -1635
rect -196 -1709 196 -1703
rect -196 -1743 -184 -1709
rect 184 -1743 196 -1709
rect -196 -1749 196 -1743
rect -252 -1793 -206 -1781
rect -252 -1969 -246 -1793
rect -212 -1969 -206 -1793
rect -252 -1981 -206 -1969
rect 206 -1793 252 -1781
rect 206 -1969 212 -1793
rect 246 -1969 252 -1793
rect 206 -1981 252 -1969
rect -196 -2019 196 -2013
rect -196 -2053 -184 -2019
rect 184 -2053 196 -2019
rect -196 -2059 196 -2053
<< properties >>
string FIXED_BBOX -343 -2138 343 2138
string gencell sky130_fd_pr__nfet_01v8_lvt
string library sky130
string parameters w 1.0 l 2.0 m 10 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
