magic
tech sky130A
magscale 1 2
timestamp 1662671833
<< error_p >>
rect -1097 930 1097 1181
rect -1097 565 1097 816
rect -1097 200 1097 451
rect -1097 -165 1097 86
rect -1097 -530 1097 -279
rect -1097 -895 1097 -644
<< nwell >>
rect -1097 930 1097 1292
rect -1097 565 1097 927
rect -1097 200 1097 562
rect -1097 -165 1097 197
rect -1097 -530 1097 -168
rect -1097 -895 1097 -533
rect -1097 -1260 1097 -898
<< pmoslvt >>
rect -1003 1030 -803 1230
rect -745 1030 -545 1230
rect -487 1030 -287 1230
rect -229 1030 -29 1230
rect 29 1030 229 1230
rect 287 1030 487 1230
rect 545 1030 745 1230
rect 803 1030 1003 1230
rect -1003 665 -803 865
rect -745 665 -545 865
rect -487 665 -287 865
rect -229 665 -29 865
rect 29 665 229 865
rect 287 665 487 865
rect 545 665 745 865
rect 803 665 1003 865
rect -1003 300 -803 500
rect -745 300 -545 500
rect -487 300 -287 500
rect -229 300 -29 500
rect 29 300 229 500
rect 287 300 487 500
rect 545 300 745 500
rect 803 300 1003 500
rect -1003 -65 -803 135
rect -745 -65 -545 135
rect -487 -65 -287 135
rect -229 -65 -29 135
rect 29 -65 229 135
rect 287 -65 487 135
rect 545 -65 745 135
rect 803 -65 1003 135
rect -1003 -430 -803 -230
rect -745 -430 -545 -230
rect -487 -430 -287 -230
rect -229 -430 -29 -230
rect 29 -430 229 -230
rect 287 -430 487 -230
rect 545 -430 745 -230
rect 803 -430 1003 -230
rect -1003 -795 -803 -595
rect -745 -795 -545 -595
rect -487 -795 -287 -595
rect -229 -795 -29 -595
rect 29 -795 229 -595
rect 287 -795 487 -595
rect 545 -795 745 -595
rect 803 -795 1003 -595
rect -1003 -1160 -803 -960
rect -745 -1160 -545 -960
rect -487 -1160 -287 -960
rect -229 -1160 -29 -960
rect 29 -1160 229 -960
rect 287 -1160 487 -960
rect 545 -1160 745 -960
rect 803 -1160 1003 -960
<< pdiff >>
rect -1061 1218 -1003 1230
rect -1061 1042 -1049 1218
rect -1015 1042 -1003 1218
rect -1061 1030 -1003 1042
rect -803 1218 -745 1230
rect -803 1042 -791 1218
rect -757 1042 -745 1218
rect -803 1030 -745 1042
rect -545 1218 -487 1230
rect -545 1042 -533 1218
rect -499 1042 -487 1218
rect -545 1030 -487 1042
rect -287 1218 -229 1230
rect -287 1042 -275 1218
rect -241 1042 -229 1218
rect -287 1030 -229 1042
rect -29 1218 29 1230
rect -29 1042 -17 1218
rect 17 1042 29 1218
rect -29 1030 29 1042
rect 229 1218 287 1230
rect 229 1042 241 1218
rect 275 1042 287 1218
rect 229 1030 287 1042
rect 487 1218 545 1230
rect 487 1042 499 1218
rect 533 1042 545 1218
rect 487 1030 545 1042
rect 745 1218 803 1230
rect 745 1042 757 1218
rect 791 1042 803 1218
rect 745 1030 803 1042
rect 1003 1218 1061 1230
rect 1003 1042 1015 1218
rect 1049 1042 1061 1218
rect 1003 1030 1061 1042
rect -1061 853 -1003 865
rect -1061 677 -1049 853
rect -1015 677 -1003 853
rect -1061 665 -1003 677
rect -803 853 -745 865
rect -803 677 -791 853
rect -757 677 -745 853
rect -803 665 -745 677
rect -545 853 -487 865
rect -545 677 -533 853
rect -499 677 -487 853
rect -545 665 -487 677
rect -287 853 -229 865
rect -287 677 -275 853
rect -241 677 -229 853
rect -287 665 -229 677
rect -29 853 29 865
rect -29 677 -17 853
rect 17 677 29 853
rect -29 665 29 677
rect 229 853 287 865
rect 229 677 241 853
rect 275 677 287 853
rect 229 665 287 677
rect 487 853 545 865
rect 487 677 499 853
rect 533 677 545 853
rect 487 665 545 677
rect 745 853 803 865
rect 745 677 757 853
rect 791 677 803 853
rect 745 665 803 677
rect 1003 853 1061 865
rect 1003 677 1015 853
rect 1049 677 1061 853
rect 1003 665 1061 677
rect -1061 488 -1003 500
rect -1061 312 -1049 488
rect -1015 312 -1003 488
rect -1061 300 -1003 312
rect -803 488 -745 500
rect -803 312 -791 488
rect -757 312 -745 488
rect -803 300 -745 312
rect -545 488 -487 500
rect -545 312 -533 488
rect -499 312 -487 488
rect -545 300 -487 312
rect -287 488 -229 500
rect -287 312 -275 488
rect -241 312 -229 488
rect -287 300 -229 312
rect -29 488 29 500
rect -29 312 -17 488
rect 17 312 29 488
rect -29 300 29 312
rect 229 488 287 500
rect 229 312 241 488
rect 275 312 287 488
rect 229 300 287 312
rect 487 488 545 500
rect 487 312 499 488
rect 533 312 545 488
rect 487 300 545 312
rect 745 488 803 500
rect 745 312 757 488
rect 791 312 803 488
rect 745 300 803 312
rect 1003 488 1061 500
rect 1003 312 1015 488
rect 1049 312 1061 488
rect 1003 300 1061 312
rect -1061 123 -1003 135
rect -1061 -53 -1049 123
rect -1015 -53 -1003 123
rect -1061 -65 -1003 -53
rect -803 123 -745 135
rect -803 -53 -791 123
rect -757 -53 -745 123
rect -803 -65 -745 -53
rect -545 123 -487 135
rect -545 -53 -533 123
rect -499 -53 -487 123
rect -545 -65 -487 -53
rect -287 123 -229 135
rect -287 -53 -275 123
rect -241 -53 -229 123
rect -287 -65 -229 -53
rect -29 123 29 135
rect -29 -53 -17 123
rect 17 -53 29 123
rect -29 -65 29 -53
rect 229 123 287 135
rect 229 -53 241 123
rect 275 -53 287 123
rect 229 -65 287 -53
rect 487 123 545 135
rect 487 -53 499 123
rect 533 -53 545 123
rect 487 -65 545 -53
rect 745 123 803 135
rect 745 -53 757 123
rect 791 -53 803 123
rect 745 -65 803 -53
rect 1003 123 1061 135
rect 1003 -53 1015 123
rect 1049 -53 1061 123
rect 1003 -65 1061 -53
rect -1061 -242 -1003 -230
rect -1061 -418 -1049 -242
rect -1015 -418 -1003 -242
rect -1061 -430 -1003 -418
rect -803 -242 -745 -230
rect -803 -418 -791 -242
rect -757 -418 -745 -242
rect -803 -430 -745 -418
rect -545 -242 -487 -230
rect -545 -418 -533 -242
rect -499 -418 -487 -242
rect -545 -430 -487 -418
rect -287 -242 -229 -230
rect -287 -418 -275 -242
rect -241 -418 -229 -242
rect -287 -430 -229 -418
rect -29 -242 29 -230
rect -29 -418 -17 -242
rect 17 -418 29 -242
rect -29 -430 29 -418
rect 229 -242 287 -230
rect 229 -418 241 -242
rect 275 -418 287 -242
rect 229 -430 287 -418
rect 487 -242 545 -230
rect 487 -418 499 -242
rect 533 -418 545 -242
rect 487 -430 545 -418
rect 745 -242 803 -230
rect 745 -418 757 -242
rect 791 -418 803 -242
rect 745 -430 803 -418
rect 1003 -242 1061 -230
rect 1003 -418 1015 -242
rect 1049 -418 1061 -242
rect 1003 -430 1061 -418
rect -1061 -607 -1003 -595
rect -1061 -783 -1049 -607
rect -1015 -783 -1003 -607
rect -1061 -795 -1003 -783
rect -803 -607 -745 -595
rect -803 -783 -791 -607
rect -757 -783 -745 -607
rect -803 -795 -745 -783
rect -545 -607 -487 -595
rect -545 -783 -533 -607
rect -499 -783 -487 -607
rect -545 -795 -487 -783
rect -287 -607 -229 -595
rect -287 -783 -275 -607
rect -241 -783 -229 -607
rect -287 -795 -229 -783
rect -29 -607 29 -595
rect -29 -783 -17 -607
rect 17 -783 29 -607
rect -29 -795 29 -783
rect 229 -607 287 -595
rect 229 -783 241 -607
rect 275 -783 287 -607
rect 229 -795 287 -783
rect 487 -607 545 -595
rect 487 -783 499 -607
rect 533 -783 545 -607
rect 487 -795 545 -783
rect 745 -607 803 -595
rect 745 -783 757 -607
rect 791 -783 803 -607
rect 745 -795 803 -783
rect 1003 -607 1061 -595
rect 1003 -783 1015 -607
rect 1049 -783 1061 -607
rect 1003 -795 1061 -783
rect -1061 -972 -1003 -960
rect -1061 -1148 -1049 -972
rect -1015 -1148 -1003 -972
rect -1061 -1160 -1003 -1148
rect -803 -972 -745 -960
rect -803 -1148 -791 -972
rect -757 -1148 -745 -972
rect -803 -1160 -745 -1148
rect -545 -972 -487 -960
rect -545 -1148 -533 -972
rect -499 -1148 -487 -972
rect -545 -1160 -487 -1148
rect -287 -972 -229 -960
rect -287 -1148 -275 -972
rect -241 -1148 -229 -972
rect -287 -1160 -229 -1148
rect -29 -972 29 -960
rect -29 -1148 -17 -972
rect 17 -1148 29 -972
rect -29 -1160 29 -1148
rect 229 -972 287 -960
rect 229 -1148 241 -972
rect 275 -1148 287 -972
rect 229 -1160 287 -1148
rect 487 -972 545 -960
rect 487 -1148 499 -972
rect 533 -1148 545 -972
rect 487 -1160 545 -1148
rect 745 -972 803 -960
rect 745 -1148 757 -972
rect 791 -1148 803 -972
rect 745 -1160 803 -1148
rect 1003 -972 1061 -960
rect 1003 -1148 1015 -972
rect 1049 -1148 1061 -972
rect 1003 -1160 1061 -1148
<< pdiffc >>
rect -1049 1042 -1015 1218
rect -791 1042 -757 1218
rect -533 1042 -499 1218
rect -275 1042 -241 1218
rect -17 1042 17 1218
rect 241 1042 275 1218
rect 499 1042 533 1218
rect 757 1042 791 1218
rect 1015 1042 1049 1218
rect -1049 677 -1015 853
rect -791 677 -757 853
rect -533 677 -499 853
rect -275 677 -241 853
rect -17 677 17 853
rect 241 677 275 853
rect 499 677 533 853
rect 757 677 791 853
rect 1015 677 1049 853
rect -1049 312 -1015 488
rect -791 312 -757 488
rect -533 312 -499 488
rect -275 312 -241 488
rect -17 312 17 488
rect 241 312 275 488
rect 499 312 533 488
rect 757 312 791 488
rect 1015 312 1049 488
rect -1049 -53 -1015 123
rect -791 -53 -757 123
rect -533 -53 -499 123
rect -275 -53 -241 123
rect -17 -53 17 123
rect 241 -53 275 123
rect 499 -53 533 123
rect 757 -53 791 123
rect 1015 -53 1049 123
rect -1049 -418 -1015 -242
rect -791 -418 -757 -242
rect -533 -418 -499 -242
rect -275 -418 -241 -242
rect -17 -418 17 -242
rect 241 -418 275 -242
rect 499 -418 533 -242
rect 757 -418 791 -242
rect 1015 -418 1049 -242
rect -1049 -783 -1015 -607
rect -791 -783 -757 -607
rect -533 -783 -499 -607
rect -275 -783 -241 -607
rect -17 -783 17 -607
rect 241 -783 275 -607
rect 499 -783 533 -607
rect 757 -783 791 -607
rect 1015 -783 1049 -607
rect -1049 -1148 -1015 -972
rect -791 -1148 -757 -972
rect -533 -1148 -499 -972
rect -275 -1148 -241 -972
rect -17 -1148 17 -972
rect 241 -1148 275 -972
rect 499 -1148 533 -972
rect 757 -1148 791 -972
rect 1015 -1148 1049 -972
<< poly >>
rect -1003 1230 -803 1256
rect -745 1230 -545 1256
rect -487 1230 -287 1256
rect -229 1230 -29 1256
rect 29 1230 229 1256
rect 287 1230 487 1256
rect 545 1230 745 1256
rect 803 1230 1003 1256
rect -1003 983 -803 1030
rect -1003 949 -987 983
rect -819 949 -803 983
rect -1003 933 -803 949
rect -745 983 -545 1030
rect -745 949 -729 983
rect -561 949 -545 983
rect -745 933 -545 949
rect -487 983 -287 1030
rect -487 949 -471 983
rect -303 949 -287 983
rect -487 933 -287 949
rect -229 983 -29 1030
rect -229 949 -213 983
rect -45 949 -29 983
rect -229 933 -29 949
rect 29 983 229 1030
rect 29 949 45 983
rect 213 949 229 983
rect 29 933 229 949
rect 287 983 487 1030
rect 287 949 303 983
rect 471 949 487 983
rect 287 933 487 949
rect 545 983 745 1030
rect 545 949 561 983
rect 729 949 745 983
rect 545 933 745 949
rect 803 983 1003 1030
rect 803 949 819 983
rect 987 949 1003 983
rect 803 933 1003 949
rect -1003 865 -803 891
rect -745 865 -545 891
rect -487 865 -287 891
rect -229 865 -29 891
rect 29 865 229 891
rect 287 865 487 891
rect 545 865 745 891
rect 803 865 1003 891
rect -1003 618 -803 665
rect -1003 584 -987 618
rect -819 584 -803 618
rect -1003 568 -803 584
rect -745 618 -545 665
rect -745 584 -729 618
rect -561 584 -545 618
rect -745 568 -545 584
rect -487 618 -287 665
rect -487 584 -471 618
rect -303 584 -287 618
rect -487 568 -287 584
rect -229 618 -29 665
rect -229 584 -213 618
rect -45 584 -29 618
rect -229 568 -29 584
rect 29 618 229 665
rect 29 584 45 618
rect 213 584 229 618
rect 29 568 229 584
rect 287 618 487 665
rect 287 584 303 618
rect 471 584 487 618
rect 287 568 487 584
rect 545 618 745 665
rect 545 584 561 618
rect 729 584 745 618
rect 545 568 745 584
rect 803 618 1003 665
rect 803 584 819 618
rect 987 584 1003 618
rect 803 568 1003 584
rect -1003 500 -803 526
rect -745 500 -545 526
rect -487 500 -287 526
rect -229 500 -29 526
rect 29 500 229 526
rect 287 500 487 526
rect 545 500 745 526
rect 803 500 1003 526
rect -1003 253 -803 300
rect -1003 219 -987 253
rect -819 219 -803 253
rect -1003 203 -803 219
rect -745 253 -545 300
rect -745 219 -729 253
rect -561 219 -545 253
rect -745 203 -545 219
rect -487 253 -287 300
rect -487 219 -471 253
rect -303 219 -287 253
rect -487 203 -287 219
rect -229 253 -29 300
rect -229 219 -213 253
rect -45 219 -29 253
rect -229 203 -29 219
rect 29 253 229 300
rect 29 219 45 253
rect 213 219 229 253
rect 29 203 229 219
rect 287 253 487 300
rect 287 219 303 253
rect 471 219 487 253
rect 287 203 487 219
rect 545 253 745 300
rect 545 219 561 253
rect 729 219 745 253
rect 545 203 745 219
rect 803 253 1003 300
rect 803 219 819 253
rect 987 219 1003 253
rect 803 203 1003 219
rect -1003 135 -803 161
rect -745 135 -545 161
rect -487 135 -287 161
rect -229 135 -29 161
rect 29 135 229 161
rect 287 135 487 161
rect 545 135 745 161
rect 803 135 1003 161
rect -1003 -112 -803 -65
rect -1003 -146 -987 -112
rect -819 -146 -803 -112
rect -1003 -162 -803 -146
rect -745 -112 -545 -65
rect -745 -146 -729 -112
rect -561 -146 -545 -112
rect -745 -162 -545 -146
rect -487 -112 -287 -65
rect -487 -146 -471 -112
rect -303 -146 -287 -112
rect -487 -162 -287 -146
rect -229 -112 -29 -65
rect -229 -146 -213 -112
rect -45 -146 -29 -112
rect -229 -162 -29 -146
rect 29 -112 229 -65
rect 29 -146 45 -112
rect 213 -146 229 -112
rect 29 -162 229 -146
rect 287 -112 487 -65
rect 287 -146 303 -112
rect 471 -146 487 -112
rect 287 -162 487 -146
rect 545 -112 745 -65
rect 545 -146 561 -112
rect 729 -146 745 -112
rect 545 -162 745 -146
rect 803 -112 1003 -65
rect 803 -146 819 -112
rect 987 -146 1003 -112
rect 803 -162 1003 -146
rect -1003 -230 -803 -204
rect -745 -230 -545 -204
rect -487 -230 -287 -204
rect -229 -230 -29 -204
rect 29 -230 229 -204
rect 287 -230 487 -204
rect 545 -230 745 -204
rect 803 -230 1003 -204
rect -1003 -477 -803 -430
rect -1003 -511 -987 -477
rect -819 -511 -803 -477
rect -1003 -527 -803 -511
rect -745 -477 -545 -430
rect -745 -511 -729 -477
rect -561 -511 -545 -477
rect -745 -527 -545 -511
rect -487 -477 -287 -430
rect -487 -511 -471 -477
rect -303 -511 -287 -477
rect -487 -527 -287 -511
rect -229 -477 -29 -430
rect -229 -511 -213 -477
rect -45 -511 -29 -477
rect -229 -527 -29 -511
rect 29 -477 229 -430
rect 29 -511 45 -477
rect 213 -511 229 -477
rect 29 -527 229 -511
rect 287 -477 487 -430
rect 287 -511 303 -477
rect 471 -511 487 -477
rect 287 -527 487 -511
rect 545 -477 745 -430
rect 545 -511 561 -477
rect 729 -511 745 -477
rect 545 -527 745 -511
rect 803 -477 1003 -430
rect 803 -511 819 -477
rect 987 -511 1003 -477
rect 803 -527 1003 -511
rect -1003 -595 -803 -569
rect -745 -595 -545 -569
rect -487 -595 -287 -569
rect -229 -595 -29 -569
rect 29 -595 229 -569
rect 287 -595 487 -569
rect 545 -595 745 -569
rect 803 -595 1003 -569
rect -1003 -842 -803 -795
rect -1003 -876 -987 -842
rect -819 -876 -803 -842
rect -1003 -892 -803 -876
rect -745 -842 -545 -795
rect -745 -876 -729 -842
rect -561 -876 -545 -842
rect -745 -892 -545 -876
rect -487 -842 -287 -795
rect -487 -876 -471 -842
rect -303 -876 -287 -842
rect -487 -892 -287 -876
rect -229 -842 -29 -795
rect -229 -876 -213 -842
rect -45 -876 -29 -842
rect -229 -892 -29 -876
rect 29 -842 229 -795
rect 29 -876 45 -842
rect 213 -876 229 -842
rect 29 -892 229 -876
rect 287 -842 487 -795
rect 287 -876 303 -842
rect 471 -876 487 -842
rect 287 -892 487 -876
rect 545 -842 745 -795
rect 545 -876 561 -842
rect 729 -876 745 -842
rect 545 -892 745 -876
rect 803 -842 1003 -795
rect 803 -876 819 -842
rect 987 -876 1003 -842
rect 803 -892 1003 -876
rect -1003 -960 -803 -934
rect -745 -960 -545 -934
rect -487 -960 -287 -934
rect -229 -960 -29 -934
rect 29 -960 229 -934
rect 287 -960 487 -934
rect 545 -960 745 -934
rect 803 -960 1003 -934
rect -1003 -1207 -803 -1160
rect -1003 -1241 -987 -1207
rect -819 -1241 -803 -1207
rect -1003 -1257 -803 -1241
rect -745 -1207 -545 -1160
rect -745 -1241 -729 -1207
rect -561 -1241 -545 -1207
rect -745 -1257 -545 -1241
rect -487 -1207 -287 -1160
rect -487 -1241 -471 -1207
rect -303 -1241 -287 -1207
rect -487 -1257 -287 -1241
rect -229 -1207 -29 -1160
rect -229 -1241 -213 -1207
rect -45 -1241 -29 -1207
rect -229 -1257 -29 -1241
rect 29 -1207 229 -1160
rect 29 -1241 45 -1207
rect 213 -1241 229 -1207
rect 29 -1257 229 -1241
rect 287 -1207 487 -1160
rect 287 -1241 303 -1207
rect 471 -1241 487 -1207
rect 287 -1257 487 -1241
rect 545 -1207 745 -1160
rect 545 -1241 561 -1207
rect 729 -1241 745 -1207
rect 545 -1257 745 -1241
rect 803 -1207 1003 -1160
rect 803 -1241 819 -1207
rect 987 -1241 1003 -1207
rect 803 -1257 1003 -1241
<< polycont >>
rect -987 949 -819 983
rect -729 949 -561 983
rect -471 949 -303 983
rect -213 949 -45 983
rect 45 949 213 983
rect 303 949 471 983
rect 561 949 729 983
rect 819 949 987 983
rect -987 584 -819 618
rect -729 584 -561 618
rect -471 584 -303 618
rect -213 584 -45 618
rect 45 584 213 618
rect 303 584 471 618
rect 561 584 729 618
rect 819 584 987 618
rect -987 219 -819 253
rect -729 219 -561 253
rect -471 219 -303 253
rect -213 219 -45 253
rect 45 219 213 253
rect 303 219 471 253
rect 561 219 729 253
rect 819 219 987 253
rect -987 -146 -819 -112
rect -729 -146 -561 -112
rect -471 -146 -303 -112
rect -213 -146 -45 -112
rect 45 -146 213 -112
rect 303 -146 471 -112
rect 561 -146 729 -112
rect 819 -146 987 -112
rect -987 -511 -819 -477
rect -729 -511 -561 -477
rect -471 -511 -303 -477
rect -213 -511 -45 -477
rect 45 -511 213 -477
rect 303 -511 471 -477
rect 561 -511 729 -477
rect 819 -511 987 -477
rect -987 -876 -819 -842
rect -729 -876 -561 -842
rect -471 -876 -303 -842
rect -213 -876 -45 -842
rect 45 -876 213 -842
rect 303 -876 471 -842
rect 561 -876 729 -842
rect 819 -876 987 -842
rect -987 -1241 -819 -1207
rect -729 -1241 -561 -1207
rect -471 -1241 -303 -1207
rect -213 -1241 -45 -1207
rect 45 -1241 213 -1207
rect 303 -1241 471 -1207
rect 561 -1241 729 -1207
rect 819 -1241 987 -1207
<< locali >>
rect -1049 1218 -1015 1234
rect -1049 1026 -1015 1042
rect -791 1218 -757 1234
rect -791 1026 -757 1042
rect -533 1218 -499 1234
rect -533 1026 -499 1042
rect -275 1218 -241 1234
rect -275 1026 -241 1042
rect -17 1218 17 1234
rect -17 1026 17 1042
rect 241 1218 275 1234
rect 241 1026 275 1042
rect 499 1218 533 1234
rect 499 1026 533 1042
rect 757 1218 791 1234
rect 757 1026 791 1042
rect 1015 1218 1049 1234
rect 1015 1026 1049 1042
rect -1003 949 -987 983
rect -819 949 -803 983
rect -745 949 -729 983
rect -561 949 -545 983
rect -487 949 -471 983
rect -303 949 -287 983
rect -229 949 -213 983
rect -45 949 -29 983
rect 29 949 45 983
rect 213 949 229 983
rect 287 949 303 983
rect 471 949 487 983
rect 545 949 561 983
rect 729 949 745 983
rect 803 949 819 983
rect 987 949 1003 983
rect -1049 853 -1015 869
rect -1049 661 -1015 677
rect -791 853 -757 869
rect -791 661 -757 677
rect -533 853 -499 869
rect -533 661 -499 677
rect -275 853 -241 869
rect -275 661 -241 677
rect -17 853 17 869
rect -17 661 17 677
rect 241 853 275 869
rect 241 661 275 677
rect 499 853 533 869
rect 499 661 533 677
rect 757 853 791 869
rect 757 661 791 677
rect 1015 853 1049 869
rect 1015 661 1049 677
rect -1003 584 -987 618
rect -819 584 -803 618
rect -745 584 -729 618
rect -561 584 -545 618
rect -487 584 -471 618
rect -303 584 -287 618
rect -229 584 -213 618
rect -45 584 -29 618
rect 29 584 45 618
rect 213 584 229 618
rect 287 584 303 618
rect 471 584 487 618
rect 545 584 561 618
rect 729 584 745 618
rect 803 584 819 618
rect 987 584 1003 618
rect -1049 488 -1015 504
rect -1049 296 -1015 312
rect -791 488 -757 504
rect -791 296 -757 312
rect -533 488 -499 504
rect -533 296 -499 312
rect -275 488 -241 504
rect -275 296 -241 312
rect -17 488 17 504
rect -17 296 17 312
rect 241 488 275 504
rect 241 296 275 312
rect 499 488 533 504
rect 499 296 533 312
rect 757 488 791 504
rect 757 296 791 312
rect 1015 488 1049 504
rect 1015 296 1049 312
rect -1003 219 -987 253
rect -819 219 -803 253
rect -745 219 -729 253
rect -561 219 -545 253
rect -487 219 -471 253
rect -303 219 -287 253
rect -229 219 -213 253
rect -45 219 -29 253
rect 29 219 45 253
rect 213 219 229 253
rect 287 219 303 253
rect 471 219 487 253
rect 545 219 561 253
rect 729 219 745 253
rect 803 219 819 253
rect 987 219 1003 253
rect -1049 123 -1015 139
rect -1049 -69 -1015 -53
rect -791 123 -757 139
rect -791 -69 -757 -53
rect -533 123 -499 139
rect -533 -69 -499 -53
rect -275 123 -241 139
rect -275 -69 -241 -53
rect -17 123 17 139
rect -17 -69 17 -53
rect 241 123 275 139
rect 241 -69 275 -53
rect 499 123 533 139
rect 499 -69 533 -53
rect 757 123 791 139
rect 757 -69 791 -53
rect 1015 123 1049 139
rect 1015 -69 1049 -53
rect -1003 -146 -987 -112
rect -819 -146 -803 -112
rect -745 -146 -729 -112
rect -561 -146 -545 -112
rect -487 -146 -471 -112
rect -303 -146 -287 -112
rect -229 -146 -213 -112
rect -45 -146 -29 -112
rect 29 -146 45 -112
rect 213 -146 229 -112
rect 287 -146 303 -112
rect 471 -146 487 -112
rect 545 -146 561 -112
rect 729 -146 745 -112
rect 803 -146 819 -112
rect 987 -146 1003 -112
rect -1049 -242 -1015 -226
rect -1049 -434 -1015 -418
rect -791 -242 -757 -226
rect -791 -434 -757 -418
rect -533 -242 -499 -226
rect -533 -434 -499 -418
rect -275 -242 -241 -226
rect -275 -434 -241 -418
rect -17 -242 17 -226
rect -17 -434 17 -418
rect 241 -242 275 -226
rect 241 -434 275 -418
rect 499 -242 533 -226
rect 499 -434 533 -418
rect 757 -242 791 -226
rect 757 -434 791 -418
rect 1015 -242 1049 -226
rect 1015 -434 1049 -418
rect -1003 -511 -987 -477
rect -819 -511 -803 -477
rect -745 -511 -729 -477
rect -561 -511 -545 -477
rect -487 -511 -471 -477
rect -303 -511 -287 -477
rect -229 -511 -213 -477
rect -45 -511 -29 -477
rect 29 -511 45 -477
rect 213 -511 229 -477
rect 287 -511 303 -477
rect 471 -511 487 -477
rect 545 -511 561 -477
rect 729 -511 745 -477
rect 803 -511 819 -477
rect 987 -511 1003 -477
rect -1049 -607 -1015 -591
rect -1049 -799 -1015 -783
rect -791 -607 -757 -591
rect -791 -799 -757 -783
rect -533 -607 -499 -591
rect -533 -799 -499 -783
rect -275 -607 -241 -591
rect -275 -799 -241 -783
rect -17 -607 17 -591
rect -17 -799 17 -783
rect 241 -607 275 -591
rect 241 -799 275 -783
rect 499 -607 533 -591
rect 499 -799 533 -783
rect 757 -607 791 -591
rect 757 -799 791 -783
rect 1015 -607 1049 -591
rect 1015 -799 1049 -783
rect -1003 -876 -987 -842
rect -819 -876 -803 -842
rect -745 -876 -729 -842
rect -561 -876 -545 -842
rect -487 -876 -471 -842
rect -303 -876 -287 -842
rect -229 -876 -213 -842
rect -45 -876 -29 -842
rect 29 -876 45 -842
rect 213 -876 229 -842
rect 287 -876 303 -842
rect 471 -876 487 -842
rect 545 -876 561 -842
rect 729 -876 745 -842
rect 803 -876 819 -842
rect 987 -876 1003 -842
rect -1049 -972 -1015 -956
rect -1049 -1164 -1015 -1148
rect -791 -972 -757 -956
rect -791 -1164 -757 -1148
rect -533 -972 -499 -956
rect -533 -1164 -499 -1148
rect -275 -972 -241 -956
rect -275 -1164 -241 -1148
rect -17 -972 17 -956
rect -17 -1164 17 -1148
rect 241 -972 275 -956
rect 241 -1164 275 -1148
rect 499 -972 533 -956
rect 499 -1164 533 -1148
rect 757 -972 791 -956
rect 757 -1164 791 -1148
rect 1015 -972 1049 -956
rect 1015 -1164 1049 -1148
rect -1003 -1241 -987 -1207
rect -819 -1241 -803 -1207
rect -745 -1241 -729 -1207
rect -561 -1241 -545 -1207
rect -487 -1241 -471 -1207
rect -303 -1241 -287 -1207
rect -229 -1241 -213 -1207
rect -45 -1241 -29 -1207
rect 29 -1241 45 -1207
rect 213 -1241 229 -1207
rect 287 -1241 303 -1207
rect 471 -1241 487 -1207
rect 545 -1241 561 -1207
rect 729 -1241 745 -1207
rect 803 -1241 819 -1207
rect 987 -1241 1003 -1207
<< viali >>
rect -1049 1042 -1015 1218
rect -791 1042 -757 1218
rect -533 1042 -499 1218
rect -275 1042 -241 1218
rect -17 1042 17 1218
rect 241 1042 275 1218
rect 499 1042 533 1218
rect 757 1042 791 1218
rect 1015 1042 1049 1218
rect -987 949 -819 983
rect -729 949 -561 983
rect -471 949 -303 983
rect -213 949 -45 983
rect 45 949 213 983
rect 303 949 471 983
rect 561 949 729 983
rect 819 949 987 983
rect -1049 677 -1015 853
rect -791 677 -757 853
rect -533 677 -499 853
rect -275 677 -241 853
rect -17 677 17 853
rect 241 677 275 853
rect 499 677 533 853
rect 757 677 791 853
rect 1015 677 1049 853
rect -987 584 -819 618
rect -729 584 -561 618
rect -471 584 -303 618
rect -213 584 -45 618
rect 45 584 213 618
rect 303 584 471 618
rect 561 584 729 618
rect 819 584 987 618
rect -1049 312 -1015 488
rect -791 312 -757 488
rect -533 312 -499 488
rect -275 312 -241 488
rect -17 312 17 488
rect 241 312 275 488
rect 499 312 533 488
rect 757 312 791 488
rect 1015 312 1049 488
rect -987 219 -819 253
rect -729 219 -561 253
rect -471 219 -303 253
rect -213 219 -45 253
rect 45 219 213 253
rect 303 219 471 253
rect 561 219 729 253
rect 819 219 987 253
rect -1049 -53 -1015 123
rect -791 -53 -757 123
rect -533 -53 -499 123
rect -275 -53 -241 123
rect -17 -53 17 123
rect 241 -53 275 123
rect 499 -53 533 123
rect 757 -53 791 123
rect 1015 -53 1049 123
rect -987 -146 -819 -112
rect -729 -146 -561 -112
rect -471 -146 -303 -112
rect -213 -146 -45 -112
rect 45 -146 213 -112
rect 303 -146 471 -112
rect 561 -146 729 -112
rect 819 -146 987 -112
rect -1049 -418 -1015 -242
rect -791 -418 -757 -242
rect -533 -418 -499 -242
rect -275 -418 -241 -242
rect -17 -418 17 -242
rect 241 -418 275 -242
rect 499 -418 533 -242
rect 757 -418 791 -242
rect 1015 -418 1049 -242
rect -987 -511 -819 -477
rect -729 -511 -561 -477
rect -471 -511 -303 -477
rect -213 -511 -45 -477
rect 45 -511 213 -477
rect 303 -511 471 -477
rect 561 -511 729 -477
rect 819 -511 987 -477
rect -1049 -783 -1015 -607
rect -791 -783 -757 -607
rect -533 -783 -499 -607
rect -275 -783 -241 -607
rect -17 -783 17 -607
rect 241 -783 275 -607
rect 499 -783 533 -607
rect 757 -783 791 -607
rect 1015 -783 1049 -607
rect -987 -876 -819 -842
rect -729 -876 -561 -842
rect -471 -876 -303 -842
rect -213 -876 -45 -842
rect 45 -876 213 -842
rect 303 -876 471 -842
rect 561 -876 729 -842
rect 819 -876 987 -842
rect -1049 -1148 -1015 -972
rect -791 -1148 -757 -972
rect -533 -1148 -499 -972
rect -275 -1148 -241 -972
rect -17 -1148 17 -972
rect 241 -1148 275 -972
rect 499 -1148 533 -972
rect 757 -1148 791 -972
rect 1015 -1148 1049 -972
rect -987 -1241 -819 -1207
rect -729 -1241 -561 -1207
rect -471 -1241 -303 -1207
rect -213 -1241 -45 -1207
rect 45 -1241 213 -1207
rect 303 -1241 471 -1207
rect 561 -1241 729 -1207
rect 819 -1241 987 -1207
<< metal1 >>
rect -1055 1218 -1009 1230
rect -1055 1042 -1049 1218
rect -1015 1042 -1009 1218
rect -1055 1030 -1009 1042
rect -797 1218 -751 1230
rect -797 1042 -791 1218
rect -757 1042 -751 1218
rect -797 1030 -751 1042
rect -539 1218 -493 1230
rect -539 1042 -533 1218
rect -499 1042 -493 1218
rect -539 1030 -493 1042
rect -281 1218 -235 1230
rect -281 1042 -275 1218
rect -241 1042 -235 1218
rect -281 1030 -235 1042
rect -23 1218 23 1230
rect -23 1042 -17 1218
rect 17 1042 23 1218
rect -23 1030 23 1042
rect 235 1218 281 1230
rect 235 1042 241 1218
rect 275 1042 281 1218
rect 235 1030 281 1042
rect 493 1218 539 1230
rect 493 1042 499 1218
rect 533 1042 539 1218
rect 493 1030 539 1042
rect 751 1218 797 1230
rect 751 1042 757 1218
rect 791 1042 797 1218
rect 751 1030 797 1042
rect 1009 1218 1055 1230
rect 1009 1042 1015 1218
rect 1049 1042 1055 1218
rect 1009 1030 1055 1042
rect -999 983 -807 989
rect -999 949 -987 983
rect -819 949 -807 983
rect -999 943 -807 949
rect -741 983 -549 989
rect -741 949 -729 983
rect -561 949 -549 983
rect -741 943 -549 949
rect -483 983 -291 989
rect -483 949 -471 983
rect -303 949 -291 983
rect -483 943 -291 949
rect -225 983 -33 989
rect -225 949 -213 983
rect -45 949 -33 983
rect -225 943 -33 949
rect 33 983 225 989
rect 33 949 45 983
rect 213 949 225 983
rect 33 943 225 949
rect 291 983 483 989
rect 291 949 303 983
rect 471 949 483 983
rect 291 943 483 949
rect 549 983 741 989
rect 549 949 561 983
rect 729 949 741 983
rect 549 943 741 949
rect 807 983 999 989
rect 807 949 819 983
rect 987 949 999 983
rect 807 943 999 949
rect -1055 853 -1009 865
rect -1055 677 -1049 853
rect -1015 677 -1009 853
rect -1055 665 -1009 677
rect -797 853 -751 865
rect -797 677 -791 853
rect -757 677 -751 853
rect -797 665 -751 677
rect -539 853 -493 865
rect -539 677 -533 853
rect -499 677 -493 853
rect -539 665 -493 677
rect -281 853 -235 865
rect -281 677 -275 853
rect -241 677 -235 853
rect -281 665 -235 677
rect -23 853 23 865
rect -23 677 -17 853
rect 17 677 23 853
rect -23 665 23 677
rect 235 853 281 865
rect 235 677 241 853
rect 275 677 281 853
rect 235 665 281 677
rect 493 853 539 865
rect 493 677 499 853
rect 533 677 539 853
rect 493 665 539 677
rect 751 853 797 865
rect 751 677 757 853
rect 791 677 797 853
rect 751 665 797 677
rect 1009 853 1055 865
rect 1009 677 1015 853
rect 1049 677 1055 853
rect 1009 665 1055 677
rect -999 618 -807 624
rect -999 584 -987 618
rect -819 584 -807 618
rect -999 578 -807 584
rect -741 618 -549 624
rect -741 584 -729 618
rect -561 584 -549 618
rect -741 578 -549 584
rect -483 618 -291 624
rect -483 584 -471 618
rect -303 584 -291 618
rect -483 578 -291 584
rect -225 618 -33 624
rect -225 584 -213 618
rect -45 584 -33 618
rect -225 578 -33 584
rect 33 618 225 624
rect 33 584 45 618
rect 213 584 225 618
rect 33 578 225 584
rect 291 618 483 624
rect 291 584 303 618
rect 471 584 483 618
rect 291 578 483 584
rect 549 618 741 624
rect 549 584 561 618
rect 729 584 741 618
rect 549 578 741 584
rect 807 618 999 624
rect 807 584 819 618
rect 987 584 999 618
rect 807 578 999 584
rect -1055 488 -1009 500
rect -1055 312 -1049 488
rect -1015 312 -1009 488
rect -1055 300 -1009 312
rect -797 488 -751 500
rect -797 312 -791 488
rect -757 312 -751 488
rect -797 300 -751 312
rect -539 488 -493 500
rect -539 312 -533 488
rect -499 312 -493 488
rect -539 300 -493 312
rect -281 488 -235 500
rect -281 312 -275 488
rect -241 312 -235 488
rect -281 300 -235 312
rect -23 488 23 500
rect -23 312 -17 488
rect 17 312 23 488
rect -23 300 23 312
rect 235 488 281 500
rect 235 312 241 488
rect 275 312 281 488
rect 235 300 281 312
rect 493 488 539 500
rect 493 312 499 488
rect 533 312 539 488
rect 493 300 539 312
rect 751 488 797 500
rect 751 312 757 488
rect 791 312 797 488
rect 751 300 797 312
rect 1009 488 1055 500
rect 1009 312 1015 488
rect 1049 312 1055 488
rect 1009 300 1055 312
rect -999 253 -807 259
rect -999 219 -987 253
rect -819 219 -807 253
rect -999 213 -807 219
rect -741 253 -549 259
rect -741 219 -729 253
rect -561 219 -549 253
rect -741 213 -549 219
rect -483 253 -291 259
rect -483 219 -471 253
rect -303 219 -291 253
rect -483 213 -291 219
rect -225 253 -33 259
rect -225 219 -213 253
rect -45 219 -33 253
rect -225 213 -33 219
rect 33 253 225 259
rect 33 219 45 253
rect 213 219 225 253
rect 33 213 225 219
rect 291 253 483 259
rect 291 219 303 253
rect 471 219 483 253
rect 291 213 483 219
rect 549 253 741 259
rect 549 219 561 253
rect 729 219 741 253
rect 549 213 741 219
rect 807 253 999 259
rect 807 219 819 253
rect 987 219 999 253
rect 807 213 999 219
rect -1055 123 -1009 135
rect -1055 -53 -1049 123
rect -1015 -53 -1009 123
rect -1055 -65 -1009 -53
rect -797 123 -751 135
rect -797 -53 -791 123
rect -757 -53 -751 123
rect -797 -65 -751 -53
rect -539 123 -493 135
rect -539 -53 -533 123
rect -499 -53 -493 123
rect -539 -65 -493 -53
rect -281 123 -235 135
rect -281 -53 -275 123
rect -241 -53 -235 123
rect -281 -65 -235 -53
rect -23 123 23 135
rect -23 -53 -17 123
rect 17 -53 23 123
rect -23 -65 23 -53
rect 235 123 281 135
rect 235 -53 241 123
rect 275 -53 281 123
rect 235 -65 281 -53
rect 493 123 539 135
rect 493 -53 499 123
rect 533 -53 539 123
rect 493 -65 539 -53
rect 751 123 797 135
rect 751 -53 757 123
rect 791 -53 797 123
rect 751 -65 797 -53
rect 1009 123 1055 135
rect 1009 -53 1015 123
rect 1049 -53 1055 123
rect 1009 -65 1055 -53
rect -999 -112 -807 -106
rect -999 -146 -987 -112
rect -819 -146 -807 -112
rect -999 -152 -807 -146
rect -741 -112 -549 -106
rect -741 -146 -729 -112
rect -561 -146 -549 -112
rect -741 -152 -549 -146
rect -483 -112 -291 -106
rect -483 -146 -471 -112
rect -303 -146 -291 -112
rect -483 -152 -291 -146
rect -225 -112 -33 -106
rect -225 -146 -213 -112
rect -45 -146 -33 -112
rect -225 -152 -33 -146
rect 33 -112 225 -106
rect 33 -146 45 -112
rect 213 -146 225 -112
rect 33 -152 225 -146
rect 291 -112 483 -106
rect 291 -146 303 -112
rect 471 -146 483 -112
rect 291 -152 483 -146
rect 549 -112 741 -106
rect 549 -146 561 -112
rect 729 -146 741 -112
rect 549 -152 741 -146
rect 807 -112 999 -106
rect 807 -146 819 -112
rect 987 -146 999 -112
rect 807 -152 999 -146
rect -1055 -242 -1009 -230
rect -1055 -418 -1049 -242
rect -1015 -418 -1009 -242
rect -1055 -430 -1009 -418
rect -797 -242 -751 -230
rect -797 -418 -791 -242
rect -757 -418 -751 -242
rect -797 -430 -751 -418
rect -539 -242 -493 -230
rect -539 -418 -533 -242
rect -499 -418 -493 -242
rect -539 -430 -493 -418
rect -281 -242 -235 -230
rect -281 -418 -275 -242
rect -241 -418 -235 -242
rect -281 -430 -235 -418
rect -23 -242 23 -230
rect -23 -418 -17 -242
rect 17 -418 23 -242
rect -23 -430 23 -418
rect 235 -242 281 -230
rect 235 -418 241 -242
rect 275 -418 281 -242
rect 235 -430 281 -418
rect 493 -242 539 -230
rect 493 -418 499 -242
rect 533 -418 539 -242
rect 493 -430 539 -418
rect 751 -242 797 -230
rect 751 -418 757 -242
rect 791 -418 797 -242
rect 751 -430 797 -418
rect 1009 -242 1055 -230
rect 1009 -418 1015 -242
rect 1049 -418 1055 -242
rect 1009 -430 1055 -418
rect -999 -477 -807 -471
rect -999 -511 -987 -477
rect -819 -511 -807 -477
rect -999 -517 -807 -511
rect -741 -477 -549 -471
rect -741 -511 -729 -477
rect -561 -511 -549 -477
rect -741 -517 -549 -511
rect -483 -477 -291 -471
rect -483 -511 -471 -477
rect -303 -511 -291 -477
rect -483 -517 -291 -511
rect -225 -477 -33 -471
rect -225 -511 -213 -477
rect -45 -511 -33 -477
rect -225 -517 -33 -511
rect 33 -477 225 -471
rect 33 -511 45 -477
rect 213 -511 225 -477
rect 33 -517 225 -511
rect 291 -477 483 -471
rect 291 -511 303 -477
rect 471 -511 483 -477
rect 291 -517 483 -511
rect 549 -477 741 -471
rect 549 -511 561 -477
rect 729 -511 741 -477
rect 549 -517 741 -511
rect 807 -477 999 -471
rect 807 -511 819 -477
rect 987 -511 999 -477
rect 807 -517 999 -511
rect -1055 -607 -1009 -595
rect -1055 -783 -1049 -607
rect -1015 -783 -1009 -607
rect -1055 -795 -1009 -783
rect -797 -607 -751 -595
rect -797 -783 -791 -607
rect -757 -783 -751 -607
rect -797 -795 -751 -783
rect -539 -607 -493 -595
rect -539 -783 -533 -607
rect -499 -783 -493 -607
rect -539 -795 -493 -783
rect -281 -607 -235 -595
rect -281 -783 -275 -607
rect -241 -783 -235 -607
rect -281 -795 -235 -783
rect -23 -607 23 -595
rect -23 -783 -17 -607
rect 17 -783 23 -607
rect -23 -795 23 -783
rect 235 -607 281 -595
rect 235 -783 241 -607
rect 275 -783 281 -607
rect 235 -795 281 -783
rect 493 -607 539 -595
rect 493 -783 499 -607
rect 533 -783 539 -607
rect 493 -795 539 -783
rect 751 -607 797 -595
rect 751 -783 757 -607
rect 791 -783 797 -607
rect 751 -795 797 -783
rect 1009 -607 1055 -595
rect 1009 -783 1015 -607
rect 1049 -783 1055 -607
rect 1009 -795 1055 -783
rect -999 -842 -807 -836
rect -999 -876 -987 -842
rect -819 -876 -807 -842
rect -999 -882 -807 -876
rect -741 -842 -549 -836
rect -741 -876 -729 -842
rect -561 -876 -549 -842
rect -741 -882 -549 -876
rect -483 -842 -291 -836
rect -483 -876 -471 -842
rect -303 -876 -291 -842
rect -483 -882 -291 -876
rect -225 -842 -33 -836
rect -225 -876 -213 -842
rect -45 -876 -33 -842
rect -225 -882 -33 -876
rect 33 -842 225 -836
rect 33 -876 45 -842
rect 213 -876 225 -842
rect 33 -882 225 -876
rect 291 -842 483 -836
rect 291 -876 303 -842
rect 471 -876 483 -842
rect 291 -882 483 -876
rect 549 -842 741 -836
rect 549 -876 561 -842
rect 729 -876 741 -842
rect 549 -882 741 -876
rect 807 -842 999 -836
rect 807 -876 819 -842
rect 987 -876 999 -842
rect 807 -882 999 -876
rect -1055 -972 -1009 -960
rect -1055 -1148 -1049 -972
rect -1015 -1148 -1009 -972
rect -1055 -1160 -1009 -1148
rect -797 -972 -751 -960
rect -797 -1148 -791 -972
rect -757 -1148 -751 -972
rect -797 -1160 -751 -1148
rect -539 -972 -493 -960
rect -539 -1148 -533 -972
rect -499 -1148 -493 -972
rect -539 -1160 -493 -1148
rect -281 -972 -235 -960
rect -281 -1148 -275 -972
rect -241 -1148 -235 -972
rect -281 -1160 -235 -1148
rect -23 -972 23 -960
rect -23 -1148 -17 -972
rect 17 -1148 23 -972
rect -23 -1160 23 -1148
rect 235 -972 281 -960
rect 235 -1148 241 -972
rect 275 -1148 281 -972
rect 235 -1160 281 -1148
rect 493 -972 539 -960
rect 493 -1148 499 -972
rect 533 -1148 539 -972
rect 493 -1160 539 -1148
rect 751 -972 797 -960
rect 751 -1148 757 -972
rect 791 -1148 797 -972
rect 751 -1160 797 -1148
rect 1009 -972 1055 -960
rect 1009 -1148 1015 -972
rect 1049 -1148 1055 -972
rect 1009 -1160 1055 -1148
rect -999 -1207 -807 -1201
rect -999 -1241 -987 -1207
rect -819 -1241 -807 -1207
rect -999 -1247 -807 -1241
rect -741 -1207 -549 -1201
rect -741 -1241 -729 -1207
rect -561 -1241 -549 -1207
rect -741 -1247 -549 -1241
rect -483 -1207 -291 -1201
rect -483 -1241 -471 -1207
rect -303 -1241 -291 -1207
rect -483 -1247 -291 -1241
rect -225 -1207 -33 -1201
rect -225 -1241 -213 -1207
rect -45 -1241 -33 -1207
rect -225 -1247 -33 -1241
rect 33 -1207 225 -1201
rect 33 -1241 45 -1207
rect 213 -1241 225 -1207
rect 33 -1247 225 -1241
rect 291 -1207 483 -1201
rect 291 -1241 303 -1207
rect 471 -1241 483 -1207
rect 291 -1247 483 -1241
rect 549 -1207 741 -1201
rect 549 -1241 561 -1207
rect 729 -1241 741 -1207
rect 549 -1247 741 -1241
rect 807 -1207 999 -1201
rect 807 -1241 819 -1207
rect 987 -1241 999 -1207
rect 807 -1247 999 -1241
<< properties >>
string gencell sky130_fd_pr__pfet_01v8_lvt
string library sky130
string parameters w 1 l 1 m 7 nf 8 diffcov 100 polycov 100 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 0 botc 1 poverlap 0 doverlap 1 lmin 0.35 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 0 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
