magic
tech sky130A
magscale 1 2
timestamp 1672344752
<< metal1 >>
rect 230 1620 240 1780
rect 320 1620 330 1780
rect 530 1620 540 1780
rect 620 1620 630 1780
rect 850 1620 860 1780
rect 940 1620 950 1780
rect 1170 1620 1180 1780
rect 1260 1620 1270 1780
rect 1490 1620 1500 1780
rect 1580 1620 1590 1780
rect 1810 1620 1820 1780
rect 1900 1620 1910 1780
rect 2110 1620 2120 1780
rect 2200 1620 2210 1780
rect 2430 1620 2440 1780
rect 2520 1620 2530 1780
rect 2750 1620 2760 1780
rect 2840 1620 2850 1780
rect 3070 1620 3080 1780
rect 3160 1620 3170 1780
rect 70 740 80 900
rect 160 740 170 900
rect 370 740 380 900
rect 460 740 470 900
rect 690 740 700 900
rect 780 740 790 900
rect 1010 740 1020 900
rect 1100 740 1110 900
rect 1330 740 1340 900
rect 1420 740 1430 900
rect 1650 740 1660 900
rect 1740 740 1750 900
rect 1950 740 1960 900
rect 2040 740 2050 900
rect 2270 740 2280 900
rect 2360 740 2370 900
rect 2590 740 2600 900
rect 2680 740 2690 900
rect 2910 740 2920 900
rect 3000 740 3010 900
rect 3230 740 3240 900
rect 3320 740 3330 900
rect 140 70 3250 130
<< via1 >>
rect 240 1620 320 1780
rect 540 1620 620 1780
rect 860 1620 940 1780
rect 1180 1620 1260 1780
rect 1500 1620 1580 1780
rect 1820 1620 1900 1780
rect 2120 1620 2200 1780
rect 2440 1620 2520 1780
rect 2760 1620 2840 1780
rect 3080 1620 3160 1780
rect 80 740 160 900
rect 380 740 460 900
rect 700 740 780 900
rect 1020 740 1100 900
rect 1340 740 1420 900
rect 1660 740 1740 900
rect 1960 740 2040 900
rect 2280 740 2360 900
rect 2600 740 2680 900
rect 2920 740 3000 900
rect 3240 740 3320 900
<< metal2 >>
rect 220 1780 3180 1800
rect 220 1620 240 1780
rect 320 1620 540 1780
rect 620 1620 860 1780
rect 940 1620 1180 1780
rect 1260 1620 1500 1780
rect 1580 1620 1820 1780
rect 1900 1620 2120 1780
rect 2200 1620 2440 1780
rect 2520 1620 2760 1780
rect 2840 1620 3080 1780
rect 3160 1620 3180 1780
rect 220 1600 3180 1620
rect 60 900 3320 920
rect 60 740 80 900
rect 160 740 380 900
rect 460 740 700 900
rect 780 740 1020 900
rect 1100 740 1340 900
rect 1420 740 1660 900
rect 1740 740 1960 900
rect 2040 740 2280 900
rect 2360 740 2600 900
rect 2680 740 2920 900
rect 3000 740 3240 900
rect 60 720 3320 740
use sky130_fd_pr__pfet_01v8_lvt_BKT746  sky130_fd_pr__pfet_01v8_lvt_BKT746_0
timestamp 1672344136
transform 1 0 1694 0 1 931
box -1747 -984 1747 984
<< end >>
