magic
tech sky130A
magscale 1 2
timestamp 1662760251
<< pwell >>
rect -307 -15948 307 15948
<< psubdiff >>
rect -271 15878 -175 15912
rect 175 15878 271 15912
rect -271 15816 -237 15878
rect 237 15816 271 15878
rect -271 -15878 -237 -15816
rect 237 -15878 271 -15816
rect -271 -15912 -175 -15878
rect 175 -15912 271 -15878
<< psubdiffcont >>
rect -175 15878 175 15912
rect -271 -15816 -237 15816
rect 237 -15816 271 15816
rect -175 -15912 175 -15878
<< xpolycontact >>
rect -141 15350 141 15782
rect -141 -15782 141 -15350
<< ppolyres >>
rect -141 -15350 141 15350
<< locali >>
rect -271 15878 -175 15912
rect 175 15878 271 15912
rect -271 15816 -237 15878
rect 237 15816 271 15878
rect -271 -15878 -237 -15816
rect 237 -15878 271 -15816
rect -271 -15912 -175 -15878
rect 175 -15912 271 -15878
<< viali >>
rect -125 15367 125 15764
rect -125 -15764 125 -15367
<< metal1 >>
rect -131 15764 131 15776
rect -131 15367 -125 15764
rect 125 15367 131 15764
rect -131 15355 131 15367
rect -131 -15367 131 -15355
rect -131 -15764 -125 -15367
rect 125 -15764 131 -15367
rect -131 -15776 131 -15764
<< res1p41 >>
rect -143 -15352 143 15352
<< properties >>
string FIXED_BBOX -254 -15895 254 15895
string gencell sky130_fd_pr__res_high_po_1p41
string library sky130
string parameters w 1.410 l 153.5 m 1 nx 1 wmin 1.410 lmin 0.50 rho 319.8 val 35.091k dummy 0 dw 0.0 term 194.82 sterm 0.0 caplen 0 guard 1 glc 1 grc 1 gtc 1 gbc 1 compatible {sky130_fd_pr__res_high_po_0p35  sky130_fd_pr__res_high_po_0p69 sky130_fd_pr__res_high_po_1p41  sky130_fd_pr__res_high_po_2p85 sky130_fd_pr__res_high_po_5p73} snake 0 full_metal 1 wmax 1.410 n_guard 0 hv_guard 0 vias 1 viagb 0 viagt 0 viagl 0 viagr 0
<< end >>
