magic
tech sky130A
magscale 1 2
timestamp 1671745787
<< error_p >>
rect -461 381 -403 387
rect -269 381 -211 387
rect -77 381 -19 387
rect 115 381 173 387
rect 307 381 365 387
rect -461 347 -449 381
rect -269 347 -257 381
rect -77 347 -65 381
rect 115 347 127 381
rect 307 347 319 381
rect -461 341 -403 347
rect -269 341 -211 347
rect -77 341 -19 347
rect 115 341 173 347
rect 307 341 365 347
rect -365 71 -307 77
rect -173 71 -115 77
rect 19 71 77 77
rect 211 71 269 77
rect 403 71 461 77
rect -365 37 -353 71
rect -173 37 -161 71
rect 19 37 31 71
rect 211 37 223 71
rect 403 37 415 71
rect -365 31 -307 37
rect -173 31 -115 37
rect 19 31 77 37
rect 211 31 269 37
rect 403 31 461 37
rect -365 -37 -307 -31
rect -173 -37 -115 -31
rect 19 -37 77 -31
rect 211 -37 269 -31
rect 403 -37 461 -31
rect -365 -71 -353 -37
rect -173 -71 -161 -37
rect 19 -71 31 -37
rect 211 -71 223 -37
rect 403 -71 415 -37
rect -365 -77 -307 -71
rect -173 -77 -115 -71
rect 19 -77 77 -71
rect 211 -77 269 -71
rect 403 -77 461 -71
rect -461 -347 -403 -341
rect -269 -347 -211 -341
rect -77 -347 -19 -341
rect 115 -347 173 -341
rect 307 -347 365 -341
rect -461 -381 -449 -347
rect -269 -381 -257 -347
rect -77 -381 -65 -347
rect 115 -381 127 -347
rect 307 -381 319 -347
rect -461 -387 -403 -381
rect -269 -387 -211 -381
rect -77 -387 -19 -381
rect 115 -387 173 -381
rect 307 -387 365 -381
<< pwell >>
rect -647 -519 647 519
<< nmoslvt >>
rect -447 109 -417 309
rect -351 109 -321 309
rect -255 109 -225 309
rect -159 109 -129 309
rect -63 109 -33 309
rect 33 109 63 309
rect 129 109 159 309
rect 225 109 255 309
rect 321 109 351 309
rect 417 109 447 309
rect -447 -309 -417 -109
rect -351 -309 -321 -109
rect -255 -309 -225 -109
rect -159 -309 -129 -109
rect -63 -309 -33 -109
rect 33 -309 63 -109
rect 129 -309 159 -109
rect 225 -309 255 -109
rect 321 -309 351 -109
rect 417 -309 447 -109
<< ndiff >>
rect -509 297 -447 309
rect -509 121 -497 297
rect -463 121 -447 297
rect -509 109 -447 121
rect -417 297 -351 309
rect -417 121 -401 297
rect -367 121 -351 297
rect -417 109 -351 121
rect -321 297 -255 309
rect -321 121 -305 297
rect -271 121 -255 297
rect -321 109 -255 121
rect -225 297 -159 309
rect -225 121 -209 297
rect -175 121 -159 297
rect -225 109 -159 121
rect -129 297 -63 309
rect -129 121 -113 297
rect -79 121 -63 297
rect -129 109 -63 121
rect -33 297 33 309
rect -33 121 -17 297
rect 17 121 33 297
rect -33 109 33 121
rect 63 297 129 309
rect 63 121 79 297
rect 113 121 129 297
rect 63 109 129 121
rect 159 297 225 309
rect 159 121 175 297
rect 209 121 225 297
rect 159 109 225 121
rect 255 297 321 309
rect 255 121 271 297
rect 305 121 321 297
rect 255 109 321 121
rect 351 297 417 309
rect 351 121 367 297
rect 401 121 417 297
rect 351 109 417 121
rect 447 297 509 309
rect 447 121 463 297
rect 497 121 509 297
rect 447 109 509 121
rect -509 -121 -447 -109
rect -509 -297 -497 -121
rect -463 -297 -447 -121
rect -509 -309 -447 -297
rect -417 -121 -351 -109
rect -417 -297 -401 -121
rect -367 -297 -351 -121
rect -417 -309 -351 -297
rect -321 -121 -255 -109
rect -321 -297 -305 -121
rect -271 -297 -255 -121
rect -321 -309 -255 -297
rect -225 -121 -159 -109
rect -225 -297 -209 -121
rect -175 -297 -159 -121
rect -225 -309 -159 -297
rect -129 -121 -63 -109
rect -129 -297 -113 -121
rect -79 -297 -63 -121
rect -129 -309 -63 -297
rect -33 -121 33 -109
rect -33 -297 -17 -121
rect 17 -297 33 -121
rect -33 -309 33 -297
rect 63 -121 129 -109
rect 63 -297 79 -121
rect 113 -297 129 -121
rect 63 -309 129 -297
rect 159 -121 225 -109
rect 159 -297 175 -121
rect 209 -297 225 -121
rect 159 -309 225 -297
rect 255 -121 321 -109
rect 255 -297 271 -121
rect 305 -297 321 -121
rect 255 -309 321 -297
rect 351 -121 417 -109
rect 351 -297 367 -121
rect 401 -297 417 -121
rect 351 -309 417 -297
rect 447 -121 509 -109
rect 447 -297 463 -121
rect 497 -297 509 -121
rect 447 -309 509 -297
<< ndiffc >>
rect -497 121 -463 297
rect -401 121 -367 297
rect -305 121 -271 297
rect -209 121 -175 297
rect -113 121 -79 297
rect -17 121 17 297
rect 79 121 113 297
rect 175 121 209 297
rect 271 121 305 297
rect 367 121 401 297
rect 463 121 497 297
rect -497 -297 -463 -121
rect -401 -297 -367 -121
rect -305 -297 -271 -121
rect -209 -297 -175 -121
rect -113 -297 -79 -121
rect -17 -297 17 -121
rect 79 -297 113 -121
rect 175 -297 209 -121
rect 271 -297 305 -121
rect 367 -297 401 -121
rect 463 -297 497 -121
<< psubdiff >>
rect -611 449 -515 483
rect 515 449 611 483
rect -611 387 -577 449
rect 577 387 611 449
rect -611 -449 -577 -387
rect 577 -449 611 -387
rect -611 -483 -515 -449
rect 515 -483 611 -449
<< psubdiffcont >>
rect -515 449 515 483
rect -611 -387 -577 387
rect 577 -387 611 387
rect -515 -483 515 -449
<< poly >>
rect -465 381 -399 397
rect -465 347 -449 381
rect -415 347 -399 381
rect -465 331 -399 347
rect -273 381 -207 397
rect -273 347 -257 381
rect -223 347 -207 381
rect -447 309 -417 331
rect -351 309 -321 335
rect -273 331 -207 347
rect -81 381 -15 397
rect -81 347 -65 381
rect -31 347 -15 381
rect -255 309 -225 331
rect -159 309 -129 335
rect -81 331 -15 347
rect 111 381 177 397
rect 111 347 127 381
rect 161 347 177 381
rect -63 309 -33 331
rect 33 309 63 335
rect 111 331 177 347
rect 303 381 369 397
rect 303 347 319 381
rect 353 347 369 381
rect 129 309 159 331
rect 225 309 255 335
rect 303 331 369 347
rect 321 309 351 331
rect 417 309 447 335
rect -447 83 -417 109
rect -351 87 -321 109
rect -369 71 -303 87
rect -255 83 -225 109
rect -159 87 -129 109
rect -369 37 -353 71
rect -319 37 -303 71
rect -369 21 -303 37
rect -177 71 -111 87
rect -63 83 -33 109
rect 33 87 63 109
rect -177 37 -161 71
rect -127 37 -111 71
rect -177 21 -111 37
rect 15 71 81 87
rect 129 83 159 109
rect 225 87 255 109
rect 15 37 31 71
rect 65 37 81 71
rect 15 21 81 37
rect 207 71 273 87
rect 321 83 351 109
rect 417 87 447 109
rect 207 37 223 71
rect 257 37 273 71
rect 207 21 273 37
rect 399 71 465 87
rect 399 37 415 71
rect 449 37 465 71
rect 399 21 465 37
rect -369 -37 -303 -21
rect -369 -71 -353 -37
rect -319 -71 -303 -37
rect -447 -109 -417 -83
rect -369 -87 -303 -71
rect -177 -37 -111 -21
rect -177 -71 -161 -37
rect -127 -71 -111 -37
rect -351 -109 -321 -87
rect -255 -109 -225 -83
rect -177 -87 -111 -71
rect 15 -37 81 -21
rect 15 -71 31 -37
rect 65 -71 81 -37
rect -159 -109 -129 -87
rect -63 -109 -33 -83
rect 15 -87 81 -71
rect 207 -37 273 -21
rect 207 -71 223 -37
rect 257 -71 273 -37
rect 33 -109 63 -87
rect 129 -109 159 -83
rect 207 -87 273 -71
rect 399 -37 465 -21
rect 399 -71 415 -37
rect 449 -71 465 -37
rect 225 -109 255 -87
rect 321 -109 351 -83
rect 399 -87 465 -71
rect 417 -109 447 -87
rect -447 -331 -417 -309
rect -465 -347 -399 -331
rect -351 -335 -321 -309
rect -255 -331 -225 -309
rect -465 -381 -449 -347
rect -415 -381 -399 -347
rect -465 -397 -399 -381
rect -273 -347 -207 -331
rect -159 -335 -129 -309
rect -63 -331 -33 -309
rect -273 -381 -257 -347
rect -223 -381 -207 -347
rect -273 -397 -207 -381
rect -81 -347 -15 -331
rect 33 -335 63 -309
rect 129 -331 159 -309
rect -81 -381 -65 -347
rect -31 -381 -15 -347
rect -81 -397 -15 -381
rect 111 -347 177 -331
rect 225 -335 255 -309
rect 321 -331 351 -309
rect 111 -381 127 -347
rect 161 -381 177 -347
rect 111 -397 177 -381
rect 303 -347 369 -331
rect 417 -335 447 -309
rect 303 -381 319 -347
rect 353 -381 369 -347
rect 303 -397 369 -381
<< polycont >>
rect -449 347 -415 381
rect -257 347 -223 381
rect -65 347 -31 381
rect 127 347 161 381
rect 319 347 353 381
rect -353 37 -319 71
rect -161 37 -127 71
rect 31 37 65 71
rect 223 37 257 71
rect 415 37 449 71
rect -353 -71 -319 -37
rect -161 -71 -127 -37
rect 31 -71 65 -37
rect 223 -71 257 -37
rect 415 -71 449 -37
rect -449 -381 -415 -347
rect -257 -381 -223 -347
rect -65 -381 -31 -347
rect 127 -381 161 -347
rect 319 -381 353 -347
<< locali >>
rect -611 449 -515 483
rect 515 449 611 483
rect -611 387 -577 449
rect 577 387 611 449
rect -465 347 -449 381
rect -415 347 -399 381
rect -273 347 -257 381
rect -223 347 -207 381
rect -81 347 -65 381
rect -31 347 -15 381
rect 111 347 127 381
rect 161 347 177 381
rect 303 347 319 381
rect 353 347 369 381
rect -497 297 -463 313
rect -497 105 -463 121
rect -401 297 -367 313
rect -401 105 -367 121
rect -305 297 -271 313
rect -305 105 -271 121
rect -209 297 -175 313
rect -209 105 -175 121
rect -113 297 -79 313
rect -113 105 -79 121
rect -17 297 17 313
rect -17 105 17 121
rect 79 297 113 313
rect 79 105 113 121
rect 175 297 209 313
rect 175 105 209 121
rect 271 297 305 313
rect 271 105 305 121
rect 367 297 401 313
rect 367 105 401 121
rect 463 297 497 313
rect 463 105 497 121
rect -369 37 -353 71
rect -319 37 -303 71
rect -177 37 -161 71
rect -127 37 -111 71
rect 15 37 31 71
rect 65 37 81 71
rect 207 37 223 71
rect 257 37 273 71
rect 399 37 415 71
rect 449 37 465 71
rect -369 -71 -353 -37
rect -319 -71 -303 -37
rect -177 -71 -161 -37
rect -127 -71 -111 -37
rect 15 -71 31 -37
rect 65 -71 81 -37
rect 207 -71 223 -37
rect 257 -71 273 -37
rect 399 -71 415 -37
rect 449 -71 465 -37
rect -497 -121 -463 -105
rect -497 -313 -463 -297
rect -401 -121 -367 -105
rect -401 -313 -367 -297
rect -305 -121 -271 -105
rect -305 -313 -271 -297
rect -209 -121 -175 -105
rect -209 -313 -175 -297
rect -113 -121 -79 -105
rect -113 -313 -79 -297
rect -17 -121 17 -105
rect -17 -313 17 -297
rect 79 -121 113 -105
rect 79 -313 113 -297
rect 175 -121 209 -105
rect 175 -313 209 -297
rect 271 -121 305 -105
rect 271 -313 305 -297
rect 367 -121 401 -105
rect 367 -313 401 -297
rect 463 -121 497 -105
rect 463 -313 497 -297
rect -465 -381 -449 -347
rect -415 -381 -399 -347
rect -273 -381 -257 -347
rect -223 -381 -207 -347
rect -81 -381 -65 -347
rect -31 -381 -15 -347
rect 111 -381 127 -347
rect 161 -381 177 -347
rect 303 -381 319 -347
rect 353 -381 369 -347
rect -611 -449 -577 -387
rect 577 -449 611 -387
rect -611 -483 -515 -449
rect 515 -483 611 -449
<< viali >>
rect -449 347 -415 381
rect -257 347 -223 381
rect -65 347 -31 381
rect 127 347 161 381
rect 319 347 353 381
rect -497 121 -463 297
rect -401 121 -367 297
rect -305 121 -271 297
rect -209 121 -175 297
rect -113 121 -79 297
rect -17 121 17 297
rect 79 121 113 297
rect 175 121 209 297
rect 271 121 305 297
rect 367 121 401 297
rect 463 121 497 297
rect -353 37 -319 71
rect -161 37 -127 71
rect 31 37 65 71
rect 223 37 257 71
rect 415 37 449 71
rect -353 -71 -319 -37
rect -161 -71 -127 -37
rect 31 -71 65 -37
rect 223 -71 257 -37
rect 415 -71 449 -37
rect -497 -297 -463 -121
rect -401 -297 -367 -121
rect -305 -297 -271 -121
rect -209 -297 -175 -121
rect -113 -297 -79 -121
rect -17 -297 17 -121
rect 79 -297 113 -121
rect 175 -297 209 -121
rect 271 -297 305 -121
rect 367 -297 401 -121
rect 463 -297 497 -121
rect -449 -381 -415 -347
rect -257 -381 -223 -347
rect -65 -381 -31 -347
rect 127 -381 161 -347
rect 319 -381 353 -347
<< metal1 >>
rect -461 381 -403 387
rect -461 347 -449 381
rect -415 347 -403 381
rect -461 341 -403 347
rect -269 381 -211 387
rect -269 347 -257 381
rect -223 347 -211 381
rect -269 341 -211 347
rect -77 381 -19 387
rect -77 347 -65 381
rect -31 347 -19 381
rect -77 341 -19 347
rect 115 381 173 387
rect 115 347 127 381
rect 161 347 173 381
rect 115 341 173 347
rect 307 381 365 387
rect 307 347 319 381
rect 353 347 365 381
rect 307 341 365 347
rect -503 297 -457 309
rect -503 121 -497 297
rect -463 121 -457 297
rect -503 109 -457 121
rect -407 297 -361 309
rect -407 121 -401 297
rect -367 121 -361 297
rect -407 109 -361 121
rect -311 297 -265 309
rect -311 121 -305 297
rect -271 121 -265 297
rect -311 109 -265 121
rect -215 297 -169 309
rect -215 121 -209 297
rect -175 121 -169 297
rect -215 109 -169 121
rect -119 297 -73 309
rect -119 121 -113 297
rect -79 121 -73 297
rect -119 109 -73 121
rect -23 297 23 309
rect -23 121 -17 297
rect 17 121 23 297
rect -23 109 23 121
rect 73 297 119 309
rect 73 121 79 297
rect 113 121 119 297
rect 73 109 119 121
rect 169 297 215 309
rect 169 121 175 297
rect 209 121 215 297
rect 169 109 215 121
rect 265 297 311 309
rect 265 121 271 297
rect 305 121 311 297
rect 265 109 311 121
rect 361 297 407 309
rect 361 121 367 297
rect 401 121 407 297
rect 361 109 407 121
rect 457 297 503 309
rect 457 121 463 297
rect 497 121 503 297
rect 457 109 503 121
rect -365 71 -307 77
rect -365 37 -353 71
rect -319 37 -307 71
rect -365 31 -307 37
rect -173 71 -115 77
rect -173 37 -161 71
rect -127 37 -115 71
rect -173 31 -115 37
rect 19 71 77 77
rect 19 37 31 71
rect 65 37 77 71
rect 19 31 77 37
rect 211 71 269 77
rect 211 37 223 71
rect 257 37 269 71
rect 211 31 269 37
rect 403 71 461 77
rect 403 37 415 71
rect 449 37 461 71
rect 403 31 461 37
rect -365 -37 -307 -31
rect -365 -71 -353 -37
rect -319 -71 -307 -37
rect -365 -77 -307 -71
rect -173 -37 -115 -31
rect -173 -71 -161 -37
rect -127 -71 -115 -37
rect -173 -77 -115 -71
rect 19 -37 77 -31
rect 19 -71 31 -37
rect 65 -71 77 -37
rect 19 -77 77 -71
rect 211 -37 269 -31
rect 211 -71 223 -37
rect 257 -71 269 -37
rect 211 -77 269 -71
rect 403 -37 461 -31
rect 403 -71 415 -37
rect 449 -71 461 -37
rect 403 -77 461 -71
rect -503 -121 -457 -109
rect -503 -297 -497 -121
rect -463 -297 -457 -121
rect -503 -309 -457 -297
rect -407 -121 -361 -109
rect -407 -297 -401 -121
rect -367 -297 -361 -121
rect -407 -309 -361 -297
rect -311 -121 -265 -109
rect -311 -297 -305 -121
rect -271 -297 -265 -121
rect -311 -309 -265 -297
rect -215 -121 -169 -109
rect -215 -297 -209 -121
rect -175 -297 -169 -121
rect -215 -309 -169 -297
rect -119 -121 -73 -109
rect -119 -297 -113 -121
rect -79 -297 -73 -121
rect -119 -309 -73 -297
rect -23 -121 23 -109
rect -23 -297 -17 -121
rect 17 -297 23 -121
rect -23 -309 23 -297
rect 73 -121 119 -109
rect 73 -297 79 -121
rect 113 -297 119 -121
rect 73 -309 119 -297
rect 169 -121 215 -109
rect 169 -297 175 -121
rect 209 -297 215 -121
rect 169 -309 215 -297
rect 265 -121 311 -109
rect 265 -297 271 -121
rect 305 -297 311 -121
rect 265 -309 311 -297
rect 361 -121 407 -109
rect 361 -297 367 -121
rect 401 -297 407 -121
rect 361 -309 407 -297
rect 457 -121 503 -109
rect 457 -297 463 -121
rect 497 -297 503 -121
rect 457 -309 503 -297
rect -461 -347 -403 -341
rect -461 -381 -449 -347
rect -415 -381 -403 -347
rect -461 -387 -403 -381
rect -269 -347 -211 -341
rect -269 -381 -257 -347
rect -223 -381 -211 -347
rect -269 -387 -211 -381
rect -77 -347 -19 -341
rect -77 -381 -65 -347
rect -31 -381 -19 -347
rect -77 -387 -19 -381
rect 115 -347 173 -341
rect 115 -381 127 -347
rect 161 -381 173 -347
rect 115 -387 173 -381
rect 307 -347 365 -341
rect 307 -381 319 -347
rect 353 -381 365 -347
rect 307 -387 365 -381
<< properties >>
string FIXED_BBOX -594 -466 594 466
string gencell sky130_fd_pr__nfet_01v8_lvt
string library sky130
string parameters w 1.0 l 0.15 m 2 nf 10 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
