magic
tech sky130A
magscale 1 2
timestamp 1671746242
<< metal3 >>
rect -750 -900 749 900
<< mimcap >>
rect -650 760 550 800
rect -650 -760 -610 760
rect 510 -760 550 760
rect -650 -800 550 -760
<< mimcapcontact >>
rect -610 -760 510 760
<< metal4 >>
rect -611 760 511 761
rect -611 -760 -610 760
rect 510 -760 511 760
rect -611 -761 511 -760
<< properties >>
string FIXED_BBOX -750 -900 650 900
string gencell sky130_fd_pr__cap_mim_m3_1
string library sky130
string parameters w 6.0 l 8.0 val 101.32 carea 2.00 cperi 0.19 nx 1 ny 1 dummy 0 square 0 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 1 tconnect 1 ccov 100
<< end >>
