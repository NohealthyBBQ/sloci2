magic
tech sky130A
magscale 1 2
timestamp 1672451792
<< locali >>
rect 11660 5680 16200 5740
rect 11660 5420 16200 5490
rect 11660 5240 16210 5290
rect 11480 4900 16380 5040
rect 11480 4100 11500 4900
rect 11600 4100 11660 4900
rect 11720 4500 13100 4660
rect 14760 4500 16140 4660
rect 11720 4220 13100 4380
rect 14760 4220 16140 4380
rect 11480 3980 11660 4100
rect 16300 4100 16380 4900
rect 16200 3980 16380 4100
rect 11480 3940 16380 3980
rect 11660 3890 16200 3940
rect 11660 3840 16210 3890
rect 11660 3590 16210 3640
rect 11670 3390 16220 3440
rect 11660 3140 16210 3190
rect 13420 1960 17060 2000
rect 12620 1000 12860 1780
rect 11100 700 12760 740
rect 11080 220 12760 280
rect 17060 -980 17220 -460
<< viali >>
rect 11500 4100 11600 4900
rect 16200 4100 16300 4900
<< metal1 >>
rect 51900 21600 52500 21800
rect 52700 21600 52710 21800
rect 33910 16220 33920 16320
rect 34020 16220 34030 16320
rect 51900 14200 52500 14400
rect 52700 14200 52710 14400
rect 11200 5700 11600 5800
rect 11200 5300 11300 5700
rect 11500 5300 11600 5700
rect 11200 4912 11600 5300
rect 16200 5700 16600 5800
rect 16200 5300 16300 5700
rect 16500 5300 16600 5700
rect 17190 5680 17200 5980
rect 17560 5680 17570 5980
rect 16200 4912 16600 5300
rect 11200 4900 11606 4912
rect 11200 4100 11500 4900
rect 11600 4100 11606 4900
rect 16194 4900 16600 4912
rect 11494 4088 11606 4100
rect 13900 4010 13970 4560
rect 16194 4100 16200 4900
rect 16300 4100 16600 4900
rect 16194 4088 16306 4100
rect 13890 3940 13900 4010
rect 13970 3940 13980 4010
rect 11530 2560 11540 2640
rect 11620 2620 11630 2640
rect 11620 2580 12440 2620
rect 11620 2560 11630 2580
rect 12220 1900 12330 2430
rect 11740 1740 12330 1900
rect 13280 2290 13370 2300
rect 13280 2220 13290 2290
rect 13360 2220 13370 2290
rect 12620 1000 12880 1780
rect 11740 800 12200 1000
rect 3000 -220 3140 140
rect 3000 -400 3020 -220
rect 3120 -400 3140 -220
rect 3000 -420 3140 -400
rect 11800 -240 11980 800
rect 13280 120 13370 2220
rect 11800 -380 11820 -240
rect 11940 -380 11980 -240
rect 11800 -420 11980 -380
rect 12700 -100 12880 80
rect 13100 20 13370 120
rect 12700 -1100 12800 -100
rect 13100 -160 13360 20
rect 16620 -100 17600 -60
rect 16620 -360 16640 -100
rect 16960 -360 17600 -100
rect 38410 -320 38420 -100
rect 38800 -320 38810 -100
rect 16620 -380 17600 -360
rect 17300 -1100 17500 -700
rect 27630 -840 27640 -620
rect 28000 -840 28010 -620
rect 38900 -1100 39100 700
rect 12590 -1300 12600 -1100
rect 12900 -1300 12910 -1100
rect 17290 -1300 17300 -1100
rect 17500 -1300 17510 -1100
rect 38890 -1300 38900 -1100
rect 39100 -1300 39110 -1100
<< via1 >>
rect 52500 21600 52700 21800
rect 33920 16220 34020 16320
rect 52500 14200 52700 14400
rect 11300 5300 11500 5700
rect 16300 5300 16500 5700
rect 17200 5680 17560 5980
rect 13900 3940 13970 4010
rect 11540 2560 11620 2640
rect 13290 2220 13360 2290
rect 3020 -400 3120 -220
rect 11820 -380 11940 -240
rect 16640 -360 16960 -100
rect 38420 -320 38800 -100
rect 27640 -840 28000 -620
rect 12600 -1300 12900 -1100
rect 17300 -1300 17500 -1100
rect 38900 -1300 39100 -1100
<< metal2 >>
rect 52500 21800 52700 21810
rect 52500 21590 52700 21600
rect 16900 21100 18800 21500
rect 19100 21400 21000 21500
rect 19100 21200 19900 21400
rect 20200 21200 21000 21400
rect 19100 21100 21000 21200
rect 21300 21400 23200 21500
rect 21300 21200 22100 21400
rect 22400 21200 23200 21400
rect 21300 21100 23200 21200
rect 23500 21400 25400 21500
rect 23500 21200 24300 21400
rect 24600 21200 25400 21400
rect 23500 21100 25400 21200
rect 25700 21400 27600 21500
rect 25700 21200 26500 21400
rect 26800 21200 27600 21400
rect 25700 21100 27600 21200
rect 27900 21400 29800 21500
rect 27900 21200 28700 21400
rect 29000 21200 29800 21400
rect 27900 21100 29800 21200
rect 30100 21400 32000 21500
rect 30100 21200 30900 21400
rect 31200 21200 32000 21400
rect 30100 21100 32000 21200
rect 32300 21400 34200 21500
rect 32300 21200 33100 21400
rect 33400 21200 34200 21400
rect 32300 21100 34200 21200
rect 17700 19880 18000 19900
rect 17700 19620 17720 19880
rect 17980 19620 18000 19880
rect 17700 19600 18000 19620
rect 33920 16320 34020 16330
rect 33920 16210 34020 16220
rect 16900 14560 34200 14900
rect 17700 14400 18000 14560
rect 17700 14190 18000 14200
rect 19900 14400 20200 14560
rect 19900 14190 20200 14200
rect 22100 14400 22400 14560
rect 22100 14190 22400 14200
rect 24300 14400 24600 14560
rect 24300 14190 24600 14200
rect 26500 14400 26800 14560
rect 26500 14190 26800 14200
rect 28700 14400 29000 14560
rect 28700 14190 29000 14200
rect 30900 14400 31200 14560
rect 30900 14190 31200 14200
rect 33100 14400 33400 14560
rect 33100 14190 33400 14200
rect 52500 14400 52700 14410
rect 52500 14190 52700 14200
rect 16660 5980 17580 6000
rect 11300 5700 11500 5710
rect 11300 5290 11500 5300
rect 16300 5700 16500 5710
rect 16300 5290 16500 5300
rect 16660 5680 17200 5980
rect 17560 5680 17580 5980
rect 16660 5660 17580 5680
rect 16660 4580 17000 5660
rect 13100 4500 13600 4520
rect 13100 4380 13120 4500
rect 13240 4380 13600 4500
rect 13100 4360 13600 4380
rect 14000 4500 14200 4510
rect 14000 4290 14200 4300
rect 16660 4220 16680 4580
rect 16980 4220 17000 4580
rect 16660 4200 17000 4220
rect 11540 4010 13980 4020
rect 11540 3940 13900 4010
rect 13970 3940 13980 4010
rect 11540 3200 11620 3940
rect 13900 3930 13970 3940
rect 7300 3000 11620 3200
rect 11540 2640 11620 3000
rect 11540 2540 11620 2560
rect 12740 2290 13370 2300
rect 12740 2220 13290 2290
rect 13360 2220 13370 2290
rect 12740 2210 13370 2220
rect 1700 1860 1800 1870
rect 1700 1750 1800 1760
rect 2160 1860 2280 1880
rect 2160 1760 2170 1860
rect 2260 1760 2280 1860
rect 1710 1660 1800 1670
rect 1710 1580 1720 1660
rect 1790 1580 1800 1660
rect 1710 1570 1800 1580
rect 2160 20 2280 1760
rect 2160 -120 2180 20
rect 2260 -120 2280 20
rect 2160 -140 2280 -120
rect 16640 -100 16960 -90
rect 3000 -220 11980 -200
rect 3000 -400 3020 -220
rect 3120 -240 11980 -220
rect 3120 -380 11820 -240
rect 11940 -380 11980 -240
rect 16640 -370 16960 -360
rect 38400 -100 38820 -80
rect 38400 -320 38420 -100
rect 38800 -320 38820 -100
rect 3120 -400 11980 -380
rect 3000 -420 11980 -400
rect 38400 -500 38820 -320
rect 27640 -620 38820 -500
rect 28000 -840 38820 -620
rect 27640 -960 38820 -840
rect 12600 -1100 12900 -1090
rect 12600 -1310 12900 -1300
rect 17300 -1100 17500 -1090
rect 17300 -1310 17500 -1300
rect 38900 -1100 39100 -1090
rect 38900 -1310 39100 -1300
<< via2 >>
rect 52500 21600 52700 21800
rect 19900 21200 20200 21400
rect 22100 21200 22400 21400
rect 24300 21200 24600 21400
rect 26500 21200 26800 21400
rect 28700 21200 29000 21400
rect 30900 21200 31200 21400
rect 33100 21200 33400 21400
rect 17720 19620 17980 19880
rect 33920 16220 34020 16320
rect 17700 14200 18000 14400
rect 19900 14200 20200 14400
rect 22100 14200 22400 14400
rect 24300 14200 24600 14400
rect 26500 14200 26800 14400
rect 28700 14200 29000 14400
rect 30900 14200 31200 14400
rect 33100 14200 33400 14400
rect 52500 14200 52700 14400
rect 11300 5300 11500 5700
rect 16300 5300 16500 5700
rect 13120 4380 13240 4500
rect 14000 4300 14200 4500
rect 16680 4220 16980 4580
rect 1700 1760 1800 1860
rect 2170 1760 2260 1860
rect 1720 1580 1790 1660
rect 2180 -120 2260 20
rect 16640 -360 16960 -100
rect 12600 -1300 12900 -1100
rect 17300 -1300 17500 -1100
rect 38900 -1300 39100 -1100
<< metal3 >>
rect 19900 21405 20200 29500
rect 22100 21405 22400 29500
rect 24300 21405 24600 29500
rect 26500 21405 26800 29500
rect 28700 21405 29000 29500
rect 30900 21405 31200 29500
rect 33100 21405 33400 29500
rect 52490 21800 52710 21805
rect 52490 21600 52500 21800
rect 52700 21600 52710 21800
rect 52490 21595 52710 21600
rect 19890 21400 20210 21405
rect 19890 21200 19900 21400
rect 20200 21200 20210 21400
rect 19890 21195 20210 21200
rect 22090 21400 22410 21405
rect 22090 21200 22100 21400
rect 22400 21200 22410 21400
rect 22090 21195 22410 21200
rect 24290 21400 24610 21405
rect 24290 21200 24300 21400
rect 24600 21200 24610 21400
rect 24290 21195 24610 21200
rect 26490 21400 26810 21405
rect 26490 21200 26500 21400
rect 26800 21200 26810 21400
rect 26490 21195 26810 21200
rect 28690 21400 29010 21405
rect 28690 21200 28700 21400
rect 29000 21200 29010 21400
rect 28690 21195 29010 21200
rect 30890 21400 31210 21405
rect 30890 21200 30900 21400
rect 31200 21200 31210 21400
rect 30890 21195 31210 21200
rect 33090 21400 33410 21405
rect 33090 21200 33100 21400
rect 33400 21200 33410 21400
rect 33090 21195 33410 21200
rect 13000 19880 18000 19900
rect 13000 19620 17720 19880
rect 17980 19620 18000 19880
rect 13000 19600 18000 19620
rect 13000 6400 13400 19600
rect 33900 16320 52100 16340
rect 33900 16220 33920 16320
rect 34020 16220 52100 16320
rect 33900 16200 52100 16220
rect 17690 14400 18010 14405
rect 17690 14200 17700 14400
rect 18000 14200 18010 14400
rect 17690 14195 18010 14200
rect 19890 14400 20210 14405
rect 19890 14200 19900 14400
rect 20200 14200 20210 14400
rect 19890 14195 20210 14200
rect 22090 14400 22410 14405
rect 22090 14200 22100 14400
rect 22400 14200 22410 14400
rect 22090 14195 22410 14200
rect 24290 14400 24610 14405
rect 24290 14200 24300 14400
rect 24600 14200 24610 14400
rect 24290 14195 24610 14200
rect 26490 14400 26810 14405
rect 26490 14200 26500 14400
rect 26800 14200 26810 14400
rect 26490 14195 26810 14200
rect 28690 14400 29010 14405
rect 28690 14200 28700 14400
rect 29000 14200 29010 14400
rect 28690 14195 29010 14200
rect 30890 14400 31210 14405
rect 30890 14200 30900 14400
rect 31200 14200 31210 14400
rect 30890 14195 31210 14200
rect 33090 14400 33410 14405
rect 33090 14200 33100 14400
rect 33400 14200 33410 14400
rect 33090 14195 33410 14200
rect 52490 14400 52710 14405
rect 52490 14200 52500 14400
rect 52700 14200 52710 14400
rect 52490 14195 52710 14200
rect 11290 5700 11510 5705
rect 11290 5300 11300 5700
rect 11500 5300 11510 5700
rect 11290 5295 11510 5300
rect 13100 4500 13260 6400
rect 16290 5700 16510 5705
rect 16290 5300 16300 5700
rect 16500 5300 16510 5700
rect 16290 5295 16510 5300
rect 13100 4380 13120 4500
rect 13240 4380 13260 4500
rect 13100 4360 13260 4380
rect 13900 4580 17000 4600
rect 13900 4500 16680 4580
rect 13900 4300 14000 4500
rect 14200 4300 16680 4500
rect 13900 4220 16680 4300
rect 16980 4220 17000 4580
rect 13900 4200 17000 4220
rect 1690 1860 2270 1870
rect 1690 1760 1700 1860
rect 1800 1760 2170 1860
rect 2260 1760 2270 1860
rect 1690 1750 2270 1760
rect 1700 1660 1810 1670
rect 1700 1580 1720 1660
rect 1790 1580 1810 1660
rect 1700 1520 1810 1580
rect 16600 40 17000 4200
rect 2160 20 17000 40
rect 2160 -120 2180 20
rect 2260 -100 17000 20
rect 2260 -120 16640 -100
rect 2160 -140 16640 -120
rect 16600 -360 16640 -140
rect 16960 -360 17000 -100
rect 16600 -400 17000 -360
rect 12590 -1100 12910 -1095
rect 12590 -1300 12600 -1100
rect 12900 -1300 12910 -1100
rect 12590 -1305 12910 -1300
rect 17290 -1100 17510 -1095
rect 17290 -1300 17300 -1100
rect 17500 -1300 17510 -1100
rect 17290 -1305 17510 -1300
rect 38890 -1100 39110 -1095
rect 38890 -1300 38900 -1100
rect 39100 -1300 39110 -1100
rect 38890 -1305 39110 -1300
<< via3 >>
rect 52500 21600 52700 21800
rect 17700 14200 18000 14400
rect 19900 14200 20200 14400
rect 22100 14200 22400 14400
rect 24300 14200 24600 14400
rect 26500 14200 26800 14400
rect 28700 14200 29000 14400
rect 30900 14200 31200 14400
rect 33100 14200 33400 14400
rect 52500 14200 52700 14400
rect 11300 5300 11500 5700
rect 16300 5300 16500 5700
rect 12600 -1300 12900 -1100
rect 17300 -1300 17500 -1100
rect 38900 -1300 39100 -1100
<< metal4 >>
rect 16600 29400 52800 29800
rect 16600 14400 16900 29400
rect 52400 21800 52800 29400
rect 52400 21600 52500 21800
rect 52700 21600 52800 21800
rect 17699 14400 18001 14401
rect 19899 14400 20201 14401
rect 22099 14400 22401 14401
rect 24299 14400 24601 14401
rect 26499 14400 26801 14401
rect 28699 14400 29001 14401
rect 30899 14400 31201 14401
rect 33099 14400 33401 14401
rect 52400 14400 52800 21600
rect 16600 14200 17700 14400
rect 18000 14200 19900 14400
rect 20200 14200 22100 14400
rect 22400 14200 24300 14400
rect 24600 14200 26500 14400
rect 26800 14200 28700 14400
rect 29000 14200 30900 14400
rect 31200 14200 33100 14400
rect 33400 14200 52500 14400
rect 52700 14200 52800 14400
rect -1400 5800 7400 6000
rect -1400 5400 -400 5800
rect 600 5400 3800 5800
rect 4800 5400 7400 5800
rect -1400 5000 7400 5400
rect -1400 3400 -800 5000
rect -1400 400 -900 3100
rect -1400 200 -800 400
rect -1400 -200 11200 200
rect -1400 -1000 -800 -200
rect 10800 -1000 11200 -200
rect 17200 -1000 17600 14200
rect 17699 14199 18001 14200
rect 19899 14199 20201 14200
rect 22099 14199 22401 14200
rect 24299 14199 24601 14200
rect 26499 14199 26801 14200
rect 28699 14199 29001 14200
rect 30899 14199 31201 14200
rect 33099 14199 33401 14200
rect 52400 -1000 52800 14200
rect -1400 -1100 52800 -1000
rect -1400 -1300 12600 -1100
rect 12900 -1300 17300 -1100
rect 17500 -1300 38900 -1100
rect 39100 -1300 52800 -1100
rect -1400 -1400 52800 -1300
<< via4 >>
rect -400 5400 600 5800
rect 3800 5400 4800 5800
rect 11200 5700 11600 5800
rect 11200 5300 11300 5700
rect 11300 5300 11500 5700
rect 11500 5300 11600 5700
rect 11200 5200 11600 5300
rect 16200 5700 16600 5800
rect 16200 5300 16300 5700
rect 16300 5300 16500 5700
rect 16500 5300 16600 5700
rect 16200 5200 16600 5300
<< metal5 >>
rect -1400 5800 17100 6000
rect -1400 5400 -400 5800
rect 600 5400 3800 5800
rect 4800 5400 11200 5800
rect -1400 5200 11200 5400
rect 11600 5200 16200 5800
rect 16600 5200 17100 5800
rect 11176 5176 11624 5200
rect 16176 5176 16624 5200
use XM_Rref  XM_Rref_0
timestamp 1662826901
transform 0 1 18173 1 0 1417
box -1417 -1173 5029 21223
use XM_current_gate  XM_current_gate_0
timestamp 1662765305
transform 1 0 11706 0 1 2648
box -106 -568 1518 462
use XM_current_gate_with_dummy  XM_current_gate_with_dummy_0
timestamp 1662842659
transform 1 0 11600 0 1 3924
box 0 -924 4660 1954
use XM_output_mirr_combined_with_dummy  XM_output_mirr_combined_with_dummy_0
timestamp 1662903677
transform 1 0 16600 0 1 14200
box -17600 -7400 35500 15000
use opamp_realcomp3_usefinger  opamp_realcomp3_usefinger_0
timestamp 1662836520
transform 1 0 4380 0 1 -594
box -5380 594 6776 6403
use sky130_fd_pr__nfet_01v8_lvt_E2U6GT  sky130_fd_pr__nfet_01v8_lvt_E2U6GT_0
timestamp 1672431769
transform 1 0 12196 0 1 1359
box -596 -679 596 679
use sky130_fd_pr__nfet_01v8_lvt_H8V8HY  sky130_fd_pr__nfet_01v8_lvt_H8V8HY_0
timestamp 1672431769
transform 1 0 13096 0 1 859
box -396 -1179 396 1179
use sky130_fd_pr__res_high_po_1p41_EL7NMZ  sky130_fd_pr__res_high_po_1p41_EL7NMZ_0
timestamp 1672432498
transform 0 -1 22598 1 0 -733
box -307 -5598 307 5598
use sky130_fd_pr__res_high_po_1p41_G3LFBQ  sky130_fd_pr__res_high_po_1p41_G3LFBQ_0
timestamp 1672432498
transform 0 1 27998 -1 0 -213
box -307 -10998 307 10998
<< labels >>
flabel metal3 13210 4940 13250 5000 0 FreeSans 960 0 0 0 C
flabel locali 14620 4940 14660 5000 0 FreeSans 960 0 0 0 C
flabel locali 13200 3850 13240 3910 0 FreeSans 960 0 0 0 C
flabel locali 14620 3870 14660 3930 0 FreeSans 960 0 0 0 C
flabel metal3 16700 2600 16900 3000 0 FreeSans 1600 0 0 0 vd4
flabel metal4 16600 21600 16900 21800 0 FreeSans 1600 0 0 0 C
flabel metal4 16600 14200 16900 14400 0 FreeSans 1600 0 0 0 C
flabel metal4 34200 14200 34500 14400 0 FreeSans 1600 0 0 0 C
flabel space 34200 21600 34500 21800 0 FreeSans 1600 0 0 0 C
flabel metal2 11020 3040 11240 3160 0 FreeSans 2400 0 0 0 Vcurrent_gate
flabel metal1 11840 100 11940 440 0 FreeSans 2400 0 0 0 Vota_bias_internal
flabel metal3 13100 6500 13300 6700 0 FreeSans 2400 0 0 0 voutb2
flabel metal3 52020 16220 52080 16320 0 FreeSans 2400 0 0 0 voutb1
flabel metal3 20000 29200 20100 29400 0 FreeSans 2400 0 0 0 Iout0
port 1 nsew
flabel metal3 22200 29200 22300 29400 0 FreeSans 2400 0 0 0 Iout1
port 2 nsew
flabel metal3 24400 29200 24500 29400 0 FreeSans 2400 0 0 0 Iout2
port 3 nsew
flabel metal3 26600 29200 26700 29400 0 FreeSans 2400 0 0 0 Iout3
port 4 nsew
flabel metal3 28800 29200 28900 29400 0 FreeSans 2400 0 0 0 Iout4
port 5 nsew
flabel metal3 31000 29200 31100 29400 0 FreeSans 2400 0 0 0 Iout5
port 6 nsew
flabel metal3 33200 29200 33300 29400 0 FreeSans 2400 0 0 0 Iout6
port 7 nsew
flabel metal3 1730 1530 1780 1550 0 FreeSans 2400 0 0 0 Vbg
port 8 nsew
flabel metal1 13300 2050 13350 2140 0 FreeSans 2400 0 0 0 Vota_bias
port 9 nsew
flabel metal5 1400 5600 2000 5800 0 FreeSans 2400 0 0 0 VDD
port 10 nsew
flabel metal4 -1200 -1000 -1000 -600 0 FreeSans 2400 0 0 0 VSS
port 11 nsew
<< end >>
