magic
tech sky130A
magscale 1 2
timestamp 1662766393
<< nmoslvt >>
rect -887 -831 -487 769
rect -429 -831 -29 769
rect 29 -831 429 769
rect 487 -831 887 769
<< ndiff >>
rect -945 757 -887 769
rect -945 -819 -933 757
rect -899 -819 -887 757
rect -945 -831 -887 -819
rect -487 757 -429 769
rect -487 -819 -475 757
rect -441 -819 -429 757
rect -487 -831 -429 -819
rect -29 757 29 769
rect -29 -819 -17 757
rect 17 -819 29 757
rect -29 -831 29 -819
rect 429 757 487 769
rect 429 -819 441 757
rect 475 -819 487 757
rect 429 -831 487 -819
rect 887 757 945 769
rect 887 -819 899 757
rect 933 -819 945 757
rect 887 -831 945 -819
<< ndiffc >>
rect -933 -819 -899 757
rect -475 -819 -441 757
rect -17 -819 17 757
rect 441 -819 475 757
rect 899 -819 933 757
<< poly >>
rect -887 841 -487 857
rect -887 807 -871 841
rect -503 807 -487 841
rect -887 769 -487 807
rect -429 841 -29 857
rect -429 807 -413 841
rect -45 807 -29 841
rect -429 769 -29 807
rect 29 841 429 857
rect 29 807 45 841
rect 413 807 429 841
rect 29 769 429 807
rect 487 841 887 857
rect 487 807 503 841
rect 871 807 887 841
rect 487 769 887 807
rect -887 -857 -487 -831
rect -429 -857 -29 -831
rect 29 -857 429 -831
rect 487 -857 887 -831
<< polycont >>
rect -871 807 -503 841
rect -413 807 -45 841
rect 45 807 413 841
rect 503 807 871 841
<< locali >>
rect -887 807 -871 841
rect -503 807 -487 841
rect -429 807 -413 841
rect -45 807 -29 841
rect 29 807 45 841
rect 413 807 429 841
rect 487 807 503 841
rect 871 807 887 841
rect -933 757 -899 773
rect -933 -835 -899 -819
rect -475 757 -441 773
rect -475 -835 -441 -819
rect -17 757 17 773
rect -17 -835 17 -819
rect 441 757 475 773
rect 441 -835 475 -819
rect 899 757 933 773
rect 899 -835 933 -819
<< viali >>
rect -871 807 -503 841
rect -413 807 -45 841
rect 45 807 413 841
rect 503 807 871 841
rect -933 -819 -899 757
rect -475 -819 -441 757
rect -17 -819 17 757
rect 441 -819 475 757
rect 899 -819 933 757
<< metal1 >>
rect -883 841 -491 847
rect -883 807 -871 841
rect -503 807 -491 841
rect -883 801 -491 807
rect -425 841 -33 847
rect -425 807 -413 841
rect -45 807 -33 841
rect -425 801 -33 807
rect 33 841 425 847
rect 33 807 45 841
rect 413 807 425 841
rect 33 801 425 807
rect 491 841 883 847
rect 491 807 503 841
rect 871 807 883 841
rect 491 801 883 807
rect -939 757 -893 769
rect -939 -819 -933 757
rect -899 -819 -893 757
rect -939 -831 -893 -819
rect -481 757 -435 769
rect -481 -819 -475 757
rect -441 -819 -435 757
rect -481 -831 -435 -819
rect -23 757 23 769
rect -23 -819 -17 757
rect 17 -819 23 757
rect -23 -831 23 -819
rect 435 757 481 769
rect 435 -819 441 757
rect 475 -819 481 757
rect 435 -831 481 -819
rect 893 757 939 769
rect 893 -819 899 757
rect 933 -819 939 757
rect 893 -831 939 -819
<< properties >>
string gencell sky130_fd_pr__nfet_01v8_lvt
string library sky130
string parameters w 8 l 2 m 1 nf 4 diffcov 100 polycov 100 guard 0 glc 0 grc 0 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 0 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 0 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
