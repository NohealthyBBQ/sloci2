magic
tech sky130A
magscale 1 2
timestamp 1662079994
<< nmos >>
rect -487 -169 -287 231
rect -229 -169 -29 231
rect 29 -169 229 231
rect 287 -169 487 231
<< ndiff >>
rect -545 219 -487 231
rect -545 -157 -533 219
rect -499 -157 -487 219
rect -545 -169 -487 -157
rect -287 219 -229 231
rect -287 -157 -275 219
rect -241 -157 -229 219
rect -287 -169 -229 -157
rect -29 219 29 231
rect -29 -157 -17 219
rect 17 -157 29 219
rect -29 -169 29 -157
rect 229 219 287 231
rect 229 -157 241 219
rect 275 -157 287 219
rect 229 -169 287 -157
rect 487 219 545 231
rect 487 -157 499 219
rect 533 -157 545 219
rect 487 -169 545 -157
<< ndiffc >>
rect -533 -157 -499 219
rect -275 -157 -241 219
rect -17 -157 17 219
rect 241 -157 275 219
rect 499 -157 533 219
<< poly >>
rect -487 231 -287 257
rect -229 231 -29 257
rect 29 231 229 257
rect 287 231 487 257
rect -487 -207 -287 -169
rect -487 -241 -471 -207
rect -303 -241 -287 -207
rect -487 -257 -287 -241
rect -229 -207 -29 -169
rect -229 -241 -213 -207
rect -45 -241 -29 -207
rect -229 -257 -29 -241
rect 29 -207 229 -169
rect 29 -241 45 -207
rect 213 -241 229 -207
rect 29 -257 229 -241
rect 287 -207 487 -169
rect 287 -241 303 -207
rect 471 -241 487 -207
rect 287 -257 487 -241
<< polycont >>
rect -471 -241 -303 -207
rect -213 -241 -45 -207
rect 45 -241 213 -207
rect 303 -241 471 -207
<< locali >>
rect -533 219 -499 235
rect -533 -173 -499 -157
rect -275 219 -241 235
rect -275 -173 -241 -157
rect -17 219 17 235
rect -17 -173 17 -157
rect 241 219 275 235
rect 241 -173 275 -157
rect 499 219 533 235
rect 499 -173 533 -157
rect -487 -241 -471 -207
rect -303 -241 -287 -207
rect -229 -241 -213 -207
rect -45 -241 -29 -207
rect 29 -241 45 -207
rect 213 -241 229 -207
rect 287 -241 303 -207
rect 471 -241 487 -207
<< viali >>
rect -533 -157 -499 219
rect -275 -157 -241 219
rect -17 -157 17 219
rect 241 -157 275 219
rect 499 -157 533 219
rect -471 -241 -303 -207
rect -213 -241 -45 -207
rect 45 -241 213 -207
rect 303 -241 471 -207
<< metal1 >>
rect -539 219 -493 231
rect -539 -157 -533 219
rect -499 -157 -493 219
rect -539 -169 -493 -157
rect -281 219 -235 231
rect -281 -157 -275 219
rect -241 -157 -235 219
rect -281 -169 -235 -157
rect -23 219 23 231
rect -23 -157 -17 219
rect 17 -157 23 219
rect -23 -169 23 -157
rect 235 219 281 231
rect 235 -157 241 219
rect 275 -157 281 219
rect 235 -169 281 -157
rect 493 219 539 231
rect 493 -157 499 219
rect 533 -157 539 219
rect 493 -169 539 -157
rect -483 -207 -291 -201
rect -483 -241 -471 -207
rect -303 -241 -291 -207
rect -483 -247 -291 -241
rect -225 -207 -33 -201
rect -225 -241 -213 -207
rect -45 -241 -33 -207
rect -225 -247 -33 -241
rect 33 -207 225 -201
rect 33 -241 45 -207
rect 213 -241 225 -207
rect 33 -247 225 -241
rect 291 -207 483 -201
rect 291 -241 303 -207
rect 471 -241 483 -207
rect 291 -247 483 -241
<< properties >>
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 2 l 1 m 1 nf 4 diffcov 100 polycov 100 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 0 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 0 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
