magic
tech sky130A
magscale 1 2
timestamp 1661907284
<< nwell >>
rect -683 -1231 683 1231
<< pmoslvt >>
rect -487 683 -287 1083
rect -229 683 -29 1083
rect 29 683 229 1083
rect 287 683 487 1083
rect -487 118 -287 518
rect -229 118 -29 518
rect 29 118 229 518
rect 287 118 487 518
rect -487 -447 -287 -47
rect -229 -447 -29 -47
rect 29 -447 229 -47
rect 287 -447 487 -47
rect -487 -1012 -287 -612
rect -229 -1012 -29 -612
rect 29 -1012 229 -612
rect 287 -1012 487 -612
<< pdiff >>
rect -545 1071 -487 1083
rect -545 695 -533 1071
rect -499 695 -487 1071
rect -545 683 -487 695
rect -287 1071 -229 1083
rect -287 695 -275 1071
rect -241 695 -229 1071
rect -287 683 -229 695
rect -29 1071 29 1083
rect -29 695 -17 1071
rect 17 695 29 1071
rect -29 683 29 695
rect 229 1071 287 1083
rect 229 695 241 1071
rect 275 695 287 1071
rect 229 683 287 695
rect 487 1071 545 1083
rect 487 695 499 1071
rect 533 695 545 1071
rect 487 683 545 695
rect -545 506 -487 518
rect -545 130 -533 506
rect -499 130 -487 506
rect -545 118 -487 130
rect -287 506 -229 518
rect -287 130 -275 506
rect -241 130 -229 506
rect -287 118 -229 130
rect -29 506 29 518
rect -29 130 -17 506
rect 17 130 29 506
rect -29 118 29 130
rect 229 506 287 518
rect 229 130 241 506
rect 275 130 287 506
rect 229 118 287 130
rect 487 506 545 518
rect 487 130 499 506
rect 533 130 545 506
rect 487 118 545 130
rect -545 -59 -487 -47
rect -545 -435 -533 -59
rect -499 -435 -487 -59
rect -545 -447 -487 -435
rect -287 -59 -229 -47
rect -287 -435 -275 -59
rect -241 -435 -229 -59
rect -287 -447 -229 -435
rect -29 -59 29 -47
rect -29 -435 -17 -59
rect 17 -435 29 -59
rect -29 -447 29 -435
rect 229 -59 287 -47
rect 229 -435 241 -59
rect 275 -435 287 -59
rect 229 -447 287 -435
rect 487 -59 545 -47
rect 487 -435 499 -59
rect 533 -435 545 -59
rect 487 -447 545 -435
rect -545 -624 -487 -612
rect -545 -1000 -533 -624
rect -499 -1000 -487 -624
rect -545 -1012 -487 -1000
rect -287 -624 -229 -612
rect -287 -1000 -275 -624
rect -241 -1000 -229 -624
rect -287 -1012 -229 -1000
rect -29 -624 29 -612
rect -29 -1000 -17 -624
rect 17 -1000 29 -624
rect -29 -1012 29 -1000
rect 229 -624 287 -612
rect 229 -1000 241 -624
rect 275 -1000 287 -624
rect 229 -1012 287 -1000
rect 487 -624 545 -612
rect 487 -1000 499 -624
rect 533 -1000 545 -624
rect 487 -1012 545 -1000
<< pdiffc >>
rect -533 695 -499 1071
rect -275 695 -241 1071
rect -17 695 17 1071
rect 241 695 275 1071
rect 499 695 533 1071
rect -533 130 -499 506
rect -275 130 -241 506
rect -17 130 17 506
rect 241 130 275 506
rect 499 130 533 506
rect -533 -435 -499 -59
rect -275 -435 -241 -59
rect -17 -435 17 -59
rect 241 -435 275 -59
rect 499 -435 533 -59
rect -533 -1000 -499 -624
rect -275 -1000 -241 -624
rect -17 -1000 17 -624
rect 241 -1000 275 -624
rect 499 -1000 533 -624
<< nsubdiff >>
rect -647 1161 -551 1195
rect 551 1161 647 1195
rect -647 1099 -613 1161
rect 613 1099 647 1161
rect -647 -1161 -613 -1099
rect 613 -1161 647 -1099
rect -647 -1195 -551 -1161
rect 551 -1195 647 -1161
<< nsubdiffcont >>
rect -551 1161 551 1195
rect -647 -1099 -613 1099
rect 613 -1099 647 1099
rect -551 -1195 551 -1161
<< poly >>
rect -487 1083 -287 1109
rect -229 1083 -29 1109
rect 29 1083 229 1109
rect 287 1083 487 1109
rect -487 636 -287 683
rect -487 602 -471 636
rect -303 602 -287 636
rect -487 586 -287 602
rect -229 636 -29 683
rect -229 602 -213 636
rect -45 602 -29 636
rect -229 586 -29 602
rect 29 636 229 683
rect 29 602 45 636
rect 213 602 229 636
rect 29 586 229 602
rect 287 636 487 683
rect 287 602 303 636
rect 471 602 487 636
rect 287 586 487 602
rect -487 518 -287 544
rect -229 518 -29 544
rect 29 518 229 544
rect 287 518 487 544
rect -487 71 -287 118
rect -487 37 -471 71
rect -303 37 -287 71
rect -487 21 -287 37
rect -229 71 -29 118
rect -229 37 -213 71
rect -45 37 -29 71
rect -229 21 -29 37
rect 29 71 229 118
rect 29 37 45 71
rect 213 37 229 71
rect 29 21 229 37
rect 287 71 487 118
rect 287 37 303 71
rect 471 37 487 71
rect 287 21 487 37
rect -487 -47 -287 -21
rect -229 -47 -29 -21
rect 29 -47 229 -21
rect 287 -47 487 -21
rect -487 -494 -287 -447
rect -487 -528 -471 -494
rect -303 -528 -287 -494
rect -487 -544 -287 -528
rect -229 -494 -29 -447
rect -229 -528 -213 -494
rect -45 -528 -29 -494
rect -229 -544 -29 -528
rect 29 -494 229 -447
rect 29 -528 45 -494
rect 213 -528 229 -494
rect 29 -544 229 -528
rect 287 -494 487 -447
rect 287 -528 303 -494
rect 471 -528 487 -494
rect 287 -544 487 -528
rect -487 -612 -287 -586
rect -229 -612 -29 -586
rect 29 -612 229 -586
rect 287 -612 487 -586
rect -487 -1059 -287 -1012
rect -487 -1093 -471 -1059
rect -303 -1093 -287 -1059
rect -487 -1109 -287 -1093
rect -229 -1059 -29 -1012
rect -229 -1093 -213 -1059
rect -45 -1093 -29 -1059
rect -229 -1109 -29 -1093
rect 29 -1059 229 -1012
rect 29 -1093 45 -1059
rect 213 -1093 229 -1059
rect 29 -1109 229 -1093
rect 287 -1059 487 -1012
rect 287 -1093 303 -1059
rect 471 -1093 487 -1059
rect 287 -1109 487 -1093
<< polycont >>
rect -471 602 -303 636
rect -213 602 -45 636
rect 45 602 213 636
rect 303 602 471 636
rect -471 37 -303 71
rect -213 37 -45 71
rect 45 37 213 71
rect 303 37 471 71
rect -471 -528 -303 -494
rect -213 -528 -45 -494
rect 45 -528 213 -494
rect 303 -528 471 -494
rect -471 -1093 -303 -1059
rect -213 -1093 -45 -1059
rect 45 -1093 213 -1059
rect 303 -1093 471 -1059
<< locali >>
rect -647 1161 -551 1195
rect 551 1161 647 1195
rect -647 1099 -613 1161
rect 613 1099 647 1161
rect -533 1071 -499 1087
rect -533 679 -499 695
rect -275 1071 -241 1087
rect -275 679 -241 695
rect -17 1071 17 1087
rect -17 679 17 695
rect 241 1071 275 1087
rect 241 679 275 695
rect 499 1071 533 1087
rect 499 679 533 695
rect -487 602 -471 636
rect -303 602 -287 636
rect -229 602 -213 636
rect -45 602 -29 636
rect 29 602 45 636
rect 213 602 229 636
rect 287 602 303 636
rect 471 602 487 636
rect -533 506 -499 522
rect -533 114 -499 130
rect -275 506 -241 522
rect -275 114 -241 130
rect -17 506 17 522
rect -17 114 17 130
rect 241 506 275 522
rect 241 114 275 130
rect 499 506 533 522
rect 499 114 533 130
rect -487 37 -471 71
rect -303 37 -287 71
rect -229 37 -213 71
rect -45 37 -29 71
rect 29 37 45 71
rect 213 37 229 71
rect 287 37 303 71
rect 471 37 487 71
rect -533 -59 -499 -43
rect -533 -451 -499 -435
rect -275 -59 -241 -43
rect -275 -451 -241 -435
rect -17 -59 17 -43
rect -17 -451 17 -435
rect 241 -59 275 -43
rect 241 -451 275 -435
rect 499 -59 533 -43
rect 499 -451 533 -435
rect -487 -528 -471 -494
rect -303 -528 -287 -494
rect -229 -528 -213 -494
rect -45 -528 -29 -494
rect 29 -528 45 -494
rect 213 -528 229 -494
rect 287 -528 303 -494
rect 471 -528 487 -494
rect -533 -624 -499 -608
rect -533 -1016 -499 -1000
rect -275 -624 -241 -608
rect -275 -1016 -241 -1000
rect -17 -624 17 -608
rect -17 -1016 17 -1000
rect 241 -624 275 -608
rect 241 -1016 275 -1000
rect 499 -624 533 -608
rect 499 -1016 533 -1000
rect -487 -1093 -471 -1059
rect -303 -1093 -287 -1059
rect -229 -1093 -213 -1059
rect -45 -1093 -29 -1059
rect 29 -1093 45 -1059
rect 213 -1093 229 -1059
rect 287 -1093 303 -1059
rect 471 -1093 487 -1059
rect -647 -1161 -613 -1099
rect 613 -1161 647 -1099
rect -647 -1195 -551 -1161
rect 551 -1195 647 -1161
<< viali >>
rect -533 695 -499 1071
rect -275 695 -241 1071
rect -17 695 17 1071
rect 241 695 275 1071
rect 499 695 533 1071
rect -471 602 -303 636
rect -213 602 -45 636
rect 45 602 213 636
rect 303 602 471 636
rect -533 130 -499 506
rect -275 130 -241 506
rect -17 130 17 506
rect 241 130 275 506
rect 499 130 533 506
rect -471 37 -303 71
rect -213 37 -45 71
rect 45 37 213 71
rect 303 37 471 71
rect -533 -435 -499 -59
rect -275 -435 -241 -59
rect -17 -435 17 -59
rect 241 -435 275 -59
rect 499 -435 533 -59
rect -471 -528 -303 -494
rect -213 -528 -45 -494
rect 45 -528 213 -494
rect 303 -528 471 -494
rect -533 -1000 -499 -624
rect -275 -1000 -241 -624
rect -17 -1000 17 -624
rect 241 -1000 275 -624
rect 499 -1000 533 -624
rect -471 -1093 -303 -1059
rect -213 -1093 -45 -1059
rect 45 -1093 213 -1059
rect 303 -1093 471 -1059
<< metal1 >>
rect -539 1071 -493 1083
rect -539 695 -533 1071
rect -499 695 -493 1071
rect -539 683 -493 695
rect -281 1071 -235 1083
rect -281 695 -275 1071
rect -241 695 -235 1071
rect -281 683 -235 695
rect -23 1071 23 1083
rect -23 695 -17 1071
rect 17 695 23 1071
rect -23 683 23 695
rect 235 1071 281 1083
rect 235 695 241 1071
rect 275 695 281 1071
rect 235 683 281 695
rect 493 1071 539 1083
rect 493 695 499 1071
rect 533 695 539 1071
rect 493 683 539 695
rect -483 636 -291 642
rect -483 602 -471 636
rect -303 602 -291 636
rect -483 596 -291 602
rect -225 636 -33 642
rect -225 602 -213 636
rect -45 602 -33 636
rect -225 596 -33 602
rect 33 636 225 642
rect 33 602 45 636
rect 213 602 225 636
rect 33 596 225 602
rect 291 636 483 642
rect 291 602 303 636
rect 471 602 483 636
rect 291 596 483 602
rect -539 506 -493 518
rect -539 130 -533 506
rect -499 130 -493 506
rect -539 118 -493 130
rect -281 506 -235 518
rect -281 130 -275 506
rect -241 130 -235 506
rect -281 118 -235 130
rect -23 506 23 518
rect -23 130 -17 506
rect 17 130 23 506
rect -23 118 23 130
rect 235 506 281 518
rect 235 130 241 506
rect 275 130 281 506
rect 235 118 281 130
rect 493 506 539 518
rect 493 130 499 506
rect 533 130 539 506
rect 493 118 539 130
rect -483 71 -291 77
rect -483 37 -471 71
rect -303 37 -291 71
rect -483 31 -291 37
rect -225 71 -33 77
rect -225 37 -213 71
rect -45 37 -33 71
rect -225 31 -33 37
rect 33 71 225 77
rect 33 37 45 71
rect 213 37 225 71
rect 33 31 225 37
rect 291 71 483 77
rect 291 37 303 71
rect 471 37 483 71
rect 291 31 483 37
rect -539 -59 -493 -47
rect -539 -435 -533 -59
rect -499 -435 -493 -59
rect -539 -447 -493 -435
rect -281 -59 -235 -47
rect -281 -435 -275 -59
rect -241 -435 -235 -59
rect -281 -447 -235 -435
rect -23 -59 23 -47
rect -23 -435 -17 -59
rect 17 -435 23 -59
rect -23 -447 23 -435
rect 235 -59 281 -47
rect 235 -435 241 -59
rect 275 -435 281 -59
rect 235 -447 281 -435
rect 493 -59 539 -47
rect 493 -435 499 -59
rect 533 -435 539 -59
rect 493 -447 539 -435
rect -483 -494 -291 -488
rect -483 -528 -471 -494
rect -303 -528 -291 -494
rect -483 -534 -291 -528
rect -225 -494 -33 -488
rect -225 -528 -213 -494
rect -45 -528 -33 -494
rect -225 -534 -33 -528
rect 33 -494 225 -488
rect 33 -528 45 -494
rect 213 -528 225 -494
rect 33 -534 225 -528
rect 291 -494 483 -488
rect 291 -528 303 -494
rect 471 -528 483 -494
rect 291 -534 483 -528
rect -539 -624 -493 -612
rect -539 -1000 -533 -624
rect -499 -1000 -493 -624
rect -539 -1012 -493 -1000
rect -281 -624 -235 -612
rect -281 -1000 -275 -624
rect -241 -1000 -235 -624
rect -281 -1012 -235 -1000
rect -23 -624 23 -612
rect -23 -1000 -17 -624
rect 17 -1000 23 -624
rect -23 -1012 23 -1000
rect 235 -624 281 -612
rect 235 -1000 241 -624
rect 275 -1000 281 -624
rect 235 -1012 281 -1000
rect 493 -624 539 -612
rect 493 -1000 499 -624
rect 533 -1000 539 -624
rect 493 -1012 539 -1000
rect -483 -1059 -291 -1053
rect -483 -1093 -471 -1059
rect -303 -1093 -291 -1059
rect -483 -1099 -291 -1093
rect -225 -1059 -33 -1053
rect -225 -1093 -213 -1059
rect -45 -1093 -33 -1059
rect -225 -1099 -33 -1093
rect 33 -1059 225 -1053
rect 33 -1093 45 -1059
rect 213 -1093 225 -1059
rect 33 -1099 225 -1093
rect 291 -1059 483 -1053
rect 291 -1093 303 -1059
rect 471 -1093 483 -1059
rect 291 -1099 483 -1093
<< properties >>
string FIXED_BBOX -630 -1178 630 1178
string gencell sky130_fd_pr__pfet_01v8_lvt
string library sky130
string parameters w 2 l 1 m 4 nf 4 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 0 botc 1 poverlap 0 doverlap 1 lmin 0.35 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
