magic
tech sky130A
magscale 1 2
timestamp 1661639644
<< pwell >>
rect -1312 -719 1312 719
<< nmoslvt >>
rect -1116 109 -716 509
rect -658 109 -258 509
rect -200 109 200 509
rect 258 109 658 509
rect 716 109 1116 509
rect -1116 -509 -716 -109
rect -658 -509 -258 -109
rect -200 -509 200 -109
rect 258 -509 658 -109
rect 716 -509 1116 -109
<< ndiff >>
rect -1174 497 -1116 509
rect -1174 121 -1162 497
rect -1128 121 -1116 497
rect -1174 109 -1116 121
rect -716 497 -658 509
rect -716 121 -704 497
rect -670 121 -658 497
rect -716 109 -658 121
rect -258 497 -200 509
rect -258 121 -246 497
rect -212 121 -200 497
rect -258 109 -200 121
rect 200 497 258 509
rect 200 121 212 497
rect 246 121 258 497
rect 200 109 258 121
rect 658 497 716 509
rect 658 121 670 497
rect 704 121 716 497
rect 658 109 716 121
rect 1116 497 1174 509
rect 1116 121 1128 497
rect 1162 121 1174 497
rect 1116 109 1174 121
rect -1174 -121 -1116 -109
rect -1174 -497 -1162 -121
rect -1128 -497 -1116 -121
rect -1174 -509 -1116 -497
rect -716 -121 -658 -109
rect -716 -497 -704 -121
rect -670 -497 -658 -121
rect -716 -509 -658 -497
rect -258 -121 -200 -109
rect -258 -497 -246 -121
rect -212 -497 -200 -121
rect -258 -509 -200 -497
rect 200 -121 258 -109
rect 200 -497 212 -121
rect 246 -497 258 -121
rect 200 -509 258 -497
rect 658 -121 716 -109
rect 658 -497 670 -121
rect 704 -497 716 -121
rect 658 -509 716 -497
rect 1116 -121 1174 -109
rect 1116 -497 1128 -121
rect 1162 -497 1174 -121
rect 1116 -509 1174 -497
<< ndiffc >>
rect -1162 121 -1128 497
rect -704 121 -670 497
rect -246 121 -212 497
rect 212 121 246 497
rect 670 121 704 497
rect 1128 121 1162 497
rect -1162 -497 -1128 -121
rect -704 -497 -670 -121
rect -246 -497 -212 -121
rect 212 -497 246 -121
rect 670 -497 704 -121
rect 1128 -497 1162 -121
<< psubdiff >>
rect -1276 649 -1180 683
rect 1180 649 1276 683
rect -1276 587 -1242 649
rect 1242 587 1276 649
rect -1276 -649 -1242 -587
rect 1242 -649 1276 -587
rect -1276 -683 -1180 -649
rect 1180 -683 1276 -649
<< psubdiffcont >>
rect -1180 649 1180 683
rect -1276 -587 -1242 587
rect 1242 -587 1276 587
rect -1180 -683 1180 -649
<< poly >>
rect -1116 581 -716 597
rect -1116 547 -1100 581
rect -732 547 -716 581
rect -1116 509 -716 547
rect -658 581 -258 597
rect -658 547 -642 581
rect -274 547 -258 581
rect -658 509 -258 547
rect -200 581 200 597
rect -200 547 -184 581
rect 184 547 200 581
rect -200 509 200 547
rect 258 581 658 597
rect 258 547 274 581
rect 642 547 658 581
rect 258 509 658 547
rect 716 581 1116 597
rect 716 547 732 581
rect 1100 547 1116 581
rect 716 509 1116 547
rect -1116 71 -716 109
rect -1116 37 -1100 71
rect -732 37 -716 71
rect -1116 21 -716 37
rect -658 71 -258 109
rect -658 37 -642 71
rect -274 37 -258 71
rect -658 21 -258 37
rect -200 71 200 109
rect -200 37 -184 71
rect 184 37 200 71
rect -200 21 200 37
rect 258 71 658 109
rect 258 37 274 71
rect 642 37 658 71
rect 258 21 658 37
rect 716 71 1116 109
rect 716 37 732 71
rect 1100 37 1116 71
rect 716 21 1116 37
rect -1116 -37 -716 -21
rect -1116 -71 -1100 -37
rect -732 -71 -716 -37
rect -1116 -109 -716 -71
rect -658 -37 -258 -21
rect -658 -71 -642 -37
rect -274 -71 -258 -37
rect -658 -109 -258 -71
rect -200 -37 200 -21
rect -200 -71 -184 -37
rect 184 -71 200 -37
rect -200 -109 200 -71
rect 258 -37 658 -21
rect 258 -71 274 -37
rect 642 -71 658 -37
rect 258 -109 658 -71
rect 716 -37 1116 -21
rect 716 -71 732 -37
rect 1100 -71 1116 -37
rect 716 -109 1116 -71
rect -1116 -547 -716 -509
rect -1116 -581 -1100 -547
rect -732 -581 -716 -547
rect -1116 -597 -716 -581
rect -658 -547 -258 -509
rect -658 -581 -642 -547
rect -274 -581 -258 -547
rect -658 -597 -258 -581
rect -200 -547 200 -509
rect -200 -581 -184 -547
rect 184 -581 200 -547
rect -200 -597 200 -581
rect 258 -547 658 -509
rect 258 -581 274 -547
rect 642 -581 658 -547
rect 258 -597 658 -581
rect 716 -547 1116 -509
rect 716 -581 732 -547
rect 1100 -581 1116 -547
rect 716 -597 1116 -581
<< polycont >>
rect -1100 547 -732 581
rect -642 547 -274 581
rect -184 547 184 581
rect 274 547 642 581
rect 732 547 1100 581
rect -1100 37 -732 71
rect -642 37 -274 71
rect -184 37 184 71
rect 274 37 642 71
rect 732 37 1100 71
rect -1100 -71 -732 -37
rect -642 -71 -274 -37
rect -184 -71 184 -37
rect 274 -71 642 -37
rect 732 -71 1100 -37
rect -1100 -581 -732 -547
rect -642 -581 -274 -547
rect -184 -581 184 -547
rect 274 -581 642 -547
rect 732 -581 1100 -547
<< locali >>
rect -1276 649 -1180 683
rect 1180 649 1276 683
rect -1276 587 -1242 649
rect 1242 587 1276 649
rect -1116 547 -1100 581
rect -732 547 -716 581
rect -658 547 -642 581
rect -274 547 -258 581
rect -200 547 -184 581
rect 184 547 200 581
rect 258 547 274 581
rect 642 547 658 581
rect 716 547 732 581
rect 1100 547 1116 581
rect -1162 497 -1128 513
rect -1162 105 -1128 121
rect -704 497 -670 513
rect -704 105 -670 121
rect -246 497 -212 513
rect -246 105 -212 121
rect 212 497 246 513
rect 212 105 246 121
rect 670 497 704 513
rect 670 105 704 121
rect 1128 497 1162 513
rect 1128 105 1162 121
rect -1116 37 -1100 71
rect -732 37 -716 71
rect -658 37 -642 71
rect -274 37 -258 71
rect -200 37 -184 71
rect 184 37 200 71
rect 258 37 274 71
rect 642 37 658 71
rect 716 37 732 71
rect 1100 37 1116 71
rect -1116 -71 -1100 -37
rect -732 -71 -716 -37
rect -658 -71 -642 -37
rect -274 -71 -258 -37
rect -200 -71 -184 -37
rect 184 -71 200 -37
rect 258 -71 274 -37
rect 642 -71 658 -37
rect 716 -71 732 -37
rect 1100 -71 1116 -37
rect -1162 -121 -1128 -105
rect -1162 -513 -1128 -497
rect -704 -121 -670 -105
rect -704 -513 -670 -497
rect -246 -121 -212 -105
rect -246 -513 -212 -497
rect 212 -121 246 -105
rect 212 -513 246 -497
rect 670 -121 704 -105
rect 670 -513 704 -497
rect 1128 -121 1162 -105
rect 1128 -513 1162 -497
rect -1116 -581 -1100 -547
rect -732 -581 -716 -547
rect -658 -581 -642 -547
rect -274 -581 -258 -547
rect -200 -581 -184 -547
rect 184 -581 200 -547
rect 258 -581 274 -547
rect 642 -581 658 -547
rect 716 -581 732 -547
rect 1100 -581 1116 -547
rect -1276 -649 -1242 -587
rect 1242 -649 1276 -587
rect -1276 -683 -1180 -649
rect 1180 -683 1276 -649
<< viali >>
rect -1100 547 -732 581
rect -642 547 -274 581
rect -184 547 184 581
rect 274 547 642 581
rect 732 547 1100 581
rect -1162 121 -1128 497
rect -704 121 -670 497
rect -246 121 -212 497
rect 212 121 246 497
rect 670 121 704 497
rect 1128 121 1162 497
rect -1100 37 -732 71
rect -642 37 -274 71
rect -184 37 184 71
rect 274 37 642 71
rect 732 37 1100 71
rect -1100 -71 -732 -37
rect -642 -71 -274 -37
rect -184 -71 184 -37
rect 274 -71 642 -37
rect 732 -71 1100 -37
rect -1162 -497 -1128 -121
rect -704 -497 -670 -121
rect -246 -497 -212 -121
rect 212 -497 246 -121
rect 670 -497 704 -121
rect 1128 -497 1162 -121
rect -1100 -581 -732 -547
rect -642 -581 -274 -547
rect -184 -581 184 -547
rect 274 -581 642 -547
rect 732 -581 1100 -547
<< metal1 >>
rect -1112 581 -720 587
rect -1112 547 -1100 581
rect -732 547 -720 581
rect -1112 541 -720 547
rect -654 581 -262 587
rect -654 547 -642 581
rect -274 547 -262 581
rect -654 541 -262 547
rect -196 581 196 587
rect -196 547 -184 581
rect 184 547 196 581
rect -196 541 196 547
rect 262 581 654 587
rect 262 547 274 581
rect 642 547 654 581
rect 262 541 654 547
rect 720 581 1112 587
rect 720 547 732 581
rect 1100 547 1112 581
rect 720 541 1112 547
rect -1168 497 -1122 509
rect -1168 121 -1162 497
rect -1128 121 -1122 497
rect -1168 109 -1122 121
rect -710 497 -664 509
rect -710 121 -704 497
rect -670 121 -664 497
rect -710 109 -664 121
rect -252 497 -206 509
rect -252 121 -246 497
rect -212 121 -206 497
rect -252 109 -206 121
rect 206 497 252 509
rect 206 121 212 497
rect 246 121 252 497
rect 206 109 252 121
rect 664 497 710 509
rect 664 121 670 497
rect 704 121 710 497
rect 664 109 710 121
rect 1122 497 1168 509
rect 1122 121 1128 497
rect 1162 121 1168 497
rect 1122 109 1168 121
rect -1112 71 -720 77
rect -1112 37 -1100 71
rect -732 37 -720 71
rect -1112 31 -720 37
rect -654 71 -262 77
rect -654 37 -642 71
rect -274 37 -262 71
rect -654 31 -262 37
rect -196 71 196 77
rect -196 37 -184 71
rect 184 37 196 71
rect -196 31 196 37
rect 262 71 654 77
rect 262 37 274 71
rect 642 37 654 71
rect 262 31 654 37
rect 720 71 1112 77
rect 720 37 732 71
rect 1100 37 1112 71
rect 720 31 1112 37
rect -1112 -37 -720 -31
rect -1112 -71 -1100 -37
rect -732 -71 -720 -37
rect -1112 -77 -720 -71
rect -654 -37 -262 -31
rect -654 -71 -642 -37
rect -274 -71 -262 -37
rect -654 -77 -262 -71
rect -196 -37 196 -31
rect -196 -71 -184 -37
rect 184 -71 196 -37
rect -196 -77 196 -71
rect 262 -37 654 -31
rect 262 -71 274 -37
rect 642 -71 654 -37
rect 262 -77 654 -71
rect 720 -37 1112 -31
rect 720 -71 732 -37
rect 1100 -71 1112 -37
rect 720 -77 1112 -71
rect -1168 -121 -1122 -109
rect -1168 -497 -1162 -121
rect -1128 -497 -1122 -121
rect -1168 -509 -1122 -497
rect -710 -121 -664 -109
rect -710 -497 -704 -121
rect -670 -497 -664 -121
rect -710 -509 -664 -497
rect -252 -121 -206 -109
rect -252 -497 -246 -121
rect -212 -497 -206 -121
rect -252 -509 -206 -497
rect 206 -121 252 -109
rect 206 -497 212 -121
rect 246 -497 252 -121
rect 206 -509 252 -497
rect 664 -121 710 -109
rect 664 -497 670 -121
rect 704 -497 710 -121
rect 664 -509 710 -497
rect 1122 -121 1168 -109
rect 1122 -497 1128 -121
rect 1162 -497 1168 -121
rect 1122 -509 1168 -497
rect -1112 -547 -720 -541
rect -1112 -581 -1100 -547
rect -732 -581 -720 -547
rect -1112 -587 -720 -581
rect -654 -547 -262 -541
rect -654 -581 -642 -547
rect -274 -581 -262 -547
rect -654 -587 -262 -581
rect -196 -547 196 -541
rect -196 -581 -184 -547
rect 184 -581 196 -547
rect -196 -587 196 -581
rect 262 -547 654 -541
rect 262 -581 274 -547
rect 642 -581 654 -547
rect 262 -587 654 -581
rect 720 -547 1112 -541
rect 720 -581 732 -547
rect 1100 -581 1112 -547
rect 720 -587 1112 -581
<< properties >>
string FIXED_BBOX -1259 -666 1259 666
string gencell sky130_fd_pr__nfet_01v8_lvt
string library sky130
string parameters w 2.0 l 2.0 m 2 nf 5 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
