magic
tech sky130A
magscale 1 2
timestamp 1672327708
<< pwell >>
rect -739 -5598 739 5598
<< psubdiff >>
rect -703 5528 -607 5562
rect 607 5528 703 5562
rect -703 -5528 -669 5528
rect 669 -5528 703 5528
rect -703 -5562 -607 -5528
rect 607 -5562 703 -5528
<< psubdiffcont >>
rect -607 5528 607 5562
rect -607 -5562 607 -5528
<< xpolycontact >>
rect -573 5000 573 5432
rect -573 -5432 573 -5000
<< xpolyres >>
rect -573 -5000 573 5000
<< locali >>
rect -703 5528 -607 5562
rect 607 5528 703 5562
rect -703 -5528 -669 5528
rect 669 -5528 703 5528
rect -703 -5562 -607 -5528
rect 607 -5562 703 -5528
<< viali >>
rect -557 5017 557 5414
rect -557 -5414 557 -5017
<< metal1 >>
rect -569 5414 569 5420
rect -569 5017 -557 5414
rect 557 5017 569 5414
rect -569 5011 569 5017
rect -569 -5017 569 -5011
rect -569 -5414 -557 -5017
rect 557 -5414 569 -5017
rect -569 -5420 569 -5414
<< res5p73 >>
rect -575 -5002 575 5002
<< properties >>
string FIXED_BBOX -686 -5545 686 5545
string gencell sky130_fd_pr__res_xhigh_po_5p73
string library sky130
string parameters w 5.73 l 50 m 1 nx 1 wmin 5.730 lmin 0.50 rho 2000 val 17.517k dummy 0 dw 0.0 term 188.2 sterm 0.0 caplen 0 wmax 5.730 guard 1 glc 0 grc 0 gtc 1 gbc 1 compatible {sky130_fd_pr__res_xhigh_po_0p35  sky130_fd_pr__res_xhigh_po_0p69 sky130_fd_pr__res_xhigh_po_1p41  sky130_fd_pr__res_xhigh_po_2p85 sky130_fd_pr__res_xhigh_po_5p73} snake 0 full_metal 1 n_guard 0 hv_guard 0 vias 1 viagb 0 viagt 0 viagl 0 viagr 0
<< end >>
