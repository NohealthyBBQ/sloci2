magic
tech sky130A
magscale 1 2
timestamp 1662733733
<< metal3 >>
rect -2450 -680 2318 680
<< mimcap >>
rect -2350 540 2250 580
rect -2350 -540 -2310 540
rect 2210 -540 2250 540
rect -2350 -580 2250 -540
<< mimcapcontact >>
rect -2310 -540 2210 540
<< metal4 >>
rect -2311 540 2211 541
rect -2311 -540 -2310 540
rect 2210 -540 2211 540
rect -2311 -541 2211 -540
<< properties >>
string FIXED_BBOX -2450 -680 2350 680
string gencell sky130_fd_pr__cap_mim_m3_1
string library sky130
string parameters w 23 l 5.8 val 277.744 carea 2.00 cperi 0.19 nx 1 ny 1 dummy 0 square 0 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 1 tconnect 1 ccov 100
<< end >>
