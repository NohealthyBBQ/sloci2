magic
tech sky130A
magscale 1 2
timestamp 1662765305
<< locali >>
rect 302 316 336 394
rect 818 316 852 394
rect 1334 316 1368 394
rect 302 -500 336 -422
rect 818 -500 852 -422
rect 1334 -500 1368 -422
<< metal1 >>
rect 30 260 40 320
rect 100 260 110 320
rect 1050 260 1060 320
rect 1120 260 1130 320
rect 530 120 540 180
rect 600 120 610 180
rect 94 27 1318 73
rect 680 -133 740 27
rect 94 -180 1318 -133
rect 530 -280 540 -220
rect 600 -280 610 -220
rect 30 -420 40 -360
rect 100 -420 110 -360
rect 1050 -420 1060 -360
rect 1120 -420 1130 -360
<< via1 >>
rect 40 260 100 320
rect 1060 260 1120 320
rect 540 120 600 180
rect 540 -280 600 -220
rect 40 -420 100 -360
rect 1060 -420 1120 -360
<< metal2 >>
rect 40 320 100 330
rect 1060 320 1120 330
rect 100 260 1060 320
rect 40 250 100 260
rect 300 -220 360 260
rect 1060 250 1120 260
rect 540 180 600 190
rect 600 120 860 180
rect 540 110 600 120
rect 540 -220 600 -210
rect 300 -280 540 -220
rect 540 -290 600 -280
rect 40 -360 100 -350
rect 800 -360 860 120
rect 1060 -360 1120 -350
rect 100 -420 1060 -360
rect 40 -430 100 -420
rect 1060 -430 1120 -420
use sky130_fd_pr__pfet_01v8_lvt_MUVY4U  sky130_fd_pr__pfet_01v8_lvt_MUVY4U_0
timestamp 1662764279
transform 1 0 706 0 1 178
box -812 -284 812 284
use sky130_fd_pr__pfet_01v8_lvt_Q24T46  sky130_fd_pr__pfet_01v8_lvt_Q24T46_0
timestamp 1662764279
transform 1 0 706 0 1 -284
box -812 -284 812 284
<< end >>
