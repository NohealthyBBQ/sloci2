magic
tech sky130A
magscale 1 2
timestamp 1662079994
<< error_p >>
rect -77 114 -19 120
rect 115 114 173 120
rect -77 80 -65 114
rect 115 80 127 114
rect -77 74 -19 80
rect 115 74 173 80
rect -173 -80 -115 -74
rect 19 -80 77 -74
rect -173 -114 -161 -80
rect 19 -114 31 -80
rect -173 -120 -115 -114
rect 19 -120 77 -114
<< nmos >>
rect -159 -42 -129 42
rect -63 -42 -33 42
rect 33 -42 63 42
rect 129 -42 159 42
<< ndiff >>
rect -221 30 -159 42
rect -221 -30 -209 30
rect -175 -30 -159 30
rect -221 -42 -159 -30
rect -129 30 -63 42
rect -129 -30 -113 30
rect -79 -30 -63 30
rect -129 -42 -63 -30
rect -33 30 33 42
rect -33 -30 -17 30
rect 17 -30 33 30
rect -33 -42 33 -30
rect 63 30 129 42
rect 63 -30 79 30
rect 113 -30 129 30
rect 63 -42 129 -30
rect 159 30 221 42
rect 159 -30 175 30
rect 209 -30 221 30
rect 159 -42 221 -30
<< ndiffc >>
rect -209 -30 -175 30
rect -113 -30 -79 30
rect -17 -30 17 30
rect 79 -30 113 30
rect 175 -30 209 30
<< poly >>
rect -81 114 -15 130
rect -81 80 -65 114
rect -31 80 -15 114
rect -159 42 -129 68
rect -81 64 -15 80
rect 111 114 177 130
rect 111 80 127 114
rect 161 80 177 114
rect -63 42 -33 64
rect 33 42 63 68
rect 111 64 177 80
rect 129 42 159 64
rect -159 -64 -129 -42
rect -177 -80 -111 -64
rect -63 -68 -33 -42
rect 33 -64 63 -42
rect -177 -114 -161 -80
rect -127 -114 -111 -80
rect -177 -130 -111 -114
rect 15 -80 81 -64
rect 129 -68 159 -42
rect 15 -114 31 -80
rect 65 -114 81 -80
rect 15 -130 81 -114
<< polycont >>
rect -65 80 -31 114
rect 127 80 161 114
rect -161 -114 -127 -80
rect 31 -114 65 -80
<< locali >>
rect -81 80 -65 114
rect -31 80 -15 114
rect 111 80 127 114
rect 161 80 177 114
rect -209 30 -175 46
rect -209 -46 -175 -30
rect -113 30 -79 46
rect -113 -46 -79 -30
rect -17 30 17 46
rect -17 -46 17 -30
rect 79 30 113 46
rect 79 -46 113 -30
rect 175 30 209 46
rect 175 -46 209 -30
rect -177 -114 -161 -80
rect -127 -114 -111 -80
rect 15 -114 31 -80
rect 65 -114 81 -80
<< viali >>
rect -65 80 -31 114
rect 127 80 161 114
rect -209 -30 -175 30
rect -113 -30 -79 30
rect -17 -30 17 30
rect 79 -30 113 30
rect 175 -30 209 30
rect -161 -114 -127 -80
rect 31 -114 65 -80
<< metal1 >>
rect -77 114 -19 120
rect -77 80 -65 114
rect -31 80 -19 114
rect -77 74 -19 80
rect 115 114 173 120
rect 115 80 127 114
rect 161 80 173 114
rect 115 74 173 80
rect -215 30 -169 42
rect -215 -30 -209 30
rect -175 -30 -169 30
rect -215 -42 -169 -30
rect -119 30 -73 42
rect -119 -30 -113 30
rect -79 -30 -73 30
rect -119 -42 -73 -30
rect -23 30 23 42
rect -23 -30 -17 30
rect 17 -30 23 30
rect -23 -42 23 -30
rect 73 30 119 42
rect 73 -30 79 30
rect 113 -30 119 30
rect 73 -42 119 -30
rect 169 30 215 42
rect 169 -30 175 30
rect 209 -30 215 30
rect 169 -42 215 -30
rect -173 -80 -115 -74
rect -173 -114 -161 -80
rect -127 -114 -115 -80
rect -173 -120 -115 -114
rect 19 -80 77 -74
rect 19 -114 31 -80
rect 65 -114 77 -80
rect 19 -120 77 -114
<< properties >>
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 0.420 l 0.150 m 1 nf 4 diffcov 100 polycov 100 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 0 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 0 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
