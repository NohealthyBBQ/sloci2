magic
tech sky130A
magscale 1 2
timestamp 1662671714
<< error_p >>
rect -968 1113 968 1364
rect -968 748 968 999
rect -968 383 968 634
rect -968 18 968 269
rect -968 -347 968 -96
rect -968 -712 968 -461
rect -968 -1077 968 -826
<< nwell >>
rect -968 1113 968 1475
rect -968 748 968 1110
rect -968 383 968 745
rect -968 18 968 380
rect -968 -347 968 15
rect -968 -712 968 -350
rect -968 -1077 968 -715
rect -968 -1442 968 -1080
<< pmoslvt >>
rect -874 1213 -674 1413
rect -616 1213 -416 1413
rect -358 1213 -158 1413
rect -100 1213 100 1413
rect 158 1213 358 1413
rect 416 1213 616 1413
rect 674 1213 874 1413
rect -874 848 -674 1048
rect -616 848 -416 1048
rect -358 848 -158 1048
rect -100 848 100 1048
rect 158 848 358 1048
rect 416 848 616 1048
rect 674 848 874 1048
rect -874 483 -674 683
rect -616 483 -416 683
rect -358 483 -158 683
rect -100 483 100 683
rect 158 483 358 683
rect 416 483 616 683
rect 674 483 874 683
rect -874 118 -674 318
rect -616 118 -416 318
rect -358 118 -158 318
rect -100 118 100 318
rect 158 118 358 318
rect 416 118 616 318
rect 674 118 874 318
rect -874 -247 -674 -47
rect -616 -247 -416 -47
rect -358 -247 -158 -47
rect -100 -247 100 -47
rect 158 -247 358 -47
rect 416 -247 616 -47
rect 674 -247 874 -47
rect -874 -612 -674 -412
rect -616 -612 -416 -412
rect -358 -612 -158 -412
rect -100 -612 100 -412
rect 158 -612 358 -412
rect 416 -612 616 -412
rect 674 -612 874 -412
rect -874 -977 -674 -777
rect -616 -977 -416 -777
rect -358 -977 -158 -777
rect -100 -977 100 -777
rect 158 -977 358 -777
rect 416 -977 616 -777
rect 674 -977 874 -777
rect -874 -1342 -674 -1142
rect -616 -1342 -416 -1142
rect -358 -1342 -158 -1142
rect -100 -1342 100 -1142
rect 158 -1342 358 -1142
rect 416 -1342 616 -1142
rect 674 -1342 874 -1142
<< pdiff >>
rect -932 1401 -874 1413
rect -932 1225 -920 1401
rect -886 1225 -874 1401
rect -932 1213 -874 1225
rect -674 1401 -616 1413
rect -674 1225 -662 1401
rect -628 1225 -616 1401
rect -674 1213 -616 1225
rect -416 1401 -358 1413
rect -416 1225 -404 1401
rect -370 1225 -358 1401
rect -416 1213 -358 1225
rect -158 1401 -100 1413
rect -158 1225 -146 1401
rect -112 1225 -100 1401
rect -158 1213 -100 1225
rect 100 1401 158 1413
rect 100 1225 112 1401
rect 146 1225 158 1401
rect 100 1213 158 1225
rect 358 1401 416 1413
rect 358 1225 370 1401
rect 404 1225 416 1401
rect 358 1213 416 1225
rect 616 1401 674 1413
rect 616 1225 628 1401
rect 662 1225 674 1401
rect 616 1213 674 1225
rect 874 1401 932 1413
rect 874 1225 886 1401
rect 920 1225 932 1401
rect 874 1213 932 1225
rect -932 1036 -874 1048
rect -932 860 -920 1036
rect -886 860 -874 1036
rect -932 848 -874 860
rect -674 1036 -616 1048
rect -674 860 -662 1036
rect -628 860 -616 1036
rect -674 848 -616 860
rect -416 1036 -358 1048
rect -416 860 -404 1036
rect -370 860 -358 1036
rect -416 848 -358 860
rect -158 1036 -100 1048
rect -158 860 -146 1036
rect -112 860 -100 1036
rect -158 848 -100 860
rect 100 1036 158 1048
rect 100 860 112 1036
rect 146 860 158 1036
rect 100 848 158 860
rect 358 1036 416 1048
rect 358 860 370 1036
rect 404 860 416 1036
rect 358 848 416 860
rect 616 1036 674 1048
rect 616 860 628 1036
rect 662 860 674 1036
rect 616 848 674 860
rect 874 1036 932 1048
rect 874 860 886 1036
rect 920 860 932 1036
rect 874 848 932 860
rect -932 671 -874 683
rect -932 495 -920 671
rect -886 495 -874 671
rect -932 483 -874 495
rect -674 671 -616 683
rect -674 495 -662 671
rect -628 495 -616 671
rect -674 483 -616 495
rect -416 671 -358 683
rect -416 495 -404 671
rect -370 495 -358 671
rect -416 483 -358 495
rect -158 671 -100 683
rect -158 495 -146 671
rect -112 495 -100 671
rect -158 483 -100 495
rect 100 671 158 683
rect 100 495 112 671
rect 146 495 158 671
rect 100 483 158 495
rect 358 671 416 683
rect 358 495 370 671
rect 404 495 416 671
rect 358 483 416 495
rect 616 671 674 683
rect 616 495 628 671
rect 662 495 674 671
rect 616 483 674 495
rect 874 671 932 683
rect 874 495 886 671
rect 920 495 932 671
rect 874 483 932 495
rect -932 306 -874 318
rect -932 130 -920 306
rect -886 130 -874 306
rect -932 118 -874 130
rect -674 306 -616 318
rect -674 130 -662 306
rect -628 130 -616 306
rect -674 118 -616 130
rect -416 306 -358 318
rect -416 130 -404 306
rect -370 130 -358 306
rect -416 118 -358 130
rect -158 306 -100 318
rect -158 130 -146 306
rect -112 130 -100 306
rect -158 118 -100 130
rect 100 306 158 318
rect 100 130 112 306
rect 146 130 158 306
rect 100 118 158 130
rect 358 306 416 318
rect 358 130 370 306
rect 404 130 416 306
rect 358 118 416 130
rect 616 306 674 318
rect 616 130 628 306
rect 662 130 674 306
rect 616 118 674 130
rect 874 306 932 318
rect 874 130 886 306
rect 920 130 932 306
rect 874 118 932 130
rect -932 -59 -874 -47
rect -932 -235 -920 -59
rect -886 -235 -874 -59
rect -932 -247 -874 -235
rect -674 -59 -616 -47
rect -674 -235 -662 -59
rect -628 -235 -616 -59
rect -674 -247 -616 -235
rect -416 -59 -358 -47
rect -416 -235 -404 -59
rect -370 -235 -358 -59
rect -416 -247 -358 -235
rect -158 -59 -100 -47
rect -158 -235 -146 -59
rect -112 -235 -100 -59
rect -158 -247 -100 -235
rect 100 -59 158 -47
rect 100 -235 112 -59
rect 146 -235 158 -59
rect 100 -247 158 -235
rect 358 -59 416 -47
rect 358 -235 370 -59
rect 404 -235 416 -59
rect 358 -247 416 -235
rect 616 -59 674 -47
rect 616 -235 628 -59
rect 662 -235 674 -59
rect 616 -247 674 -235
rect 874 -59 932 -47
rect 874 -235 886 -59
rect 920 -235 932 -59
rect 874 -247 932 -235
rect -932 -424 -874 -412
rect -932 -600 -920 -424
rect -886 -600 -874 -424
rect -932 -612 -874 -600
rect -674 -424 -616 -412
rect -674 -600 -662 -424
rect -628 -600 -616 -424
rect -674 -612 -616 -600
rect -416 -424 -358 -412
rect -416 -600 -404 -424
rect -370 -600 -358 -424
rect -416 -612 -358 -600
rect -158 -424 -100 -412
rect -158 -600 -146 -424
rect -112 -600 -100 -424
rect -158 -612 -100 -600
rect 100 -424 158 -412
rect 100 -600 112 -424
rect 146 -600 158 -424
rect 100 -612 158 -600
rect 358 -424 416 -412
rect 358 -600 370 -424
rect 404 -600 416 -424
rect 358 -612 416 -600
rect 616 -424 674 -412
rect 616 -600 628 -424
rect 662 -600 674 -424
rect 616 -612 674 -600
rect 874 -424 932 -412
rect 874 -600 886 -424
rect 920 -600 932 -424
rect 874 -612 932 -600
rect -932 -789 -874 -777
rect -932 -965 -920 -789
rect -886 -965 -874 -789
rect -932 -977 -874 -965
rect -674 -789 -616 -777
rect -674 -965 -662 -789
rect -628 -965 -616 -789
rect -674 -977 -616 -965
rect -416 -789 -358 -777
rect -416 -965 -404 -789
rect -370 -965 -358 -789
rect -416 -977 -358 -965
rect -158 -789 -100 -777
rect -158 -965 -146 -789
rect -112 -965 -100 -789
rect -158 -977 -100 -965
rect 100 -789 158 -777
rect 100 -965 112 -789
rect 146 -965 158 -789
rect 100 -977 158 -965
rect 358 -789 416 -777
rect 358 -965 370 -789
rect 404 -965 416 -789
rect 358 -977 416 -965
rect 616 -789 674 -777
rect 616 -965 628 -789
rect 662 -965 674 -789
rect 616 -977 674 -965
rect 874 -789 932 -777
rect 874 -965 886 -789
rect 920 -965 932 -789
rect 874 -977 932 -965
rect -932 -1154 -874 -1142
rect -932 -1330 -920 -1154
rect -886 -1330 -874 -1154
rect -932 -1342 -874 -1330
rect -674 -1154 -616 -1142
rect -674 -1330 -662 -1154
rect -628 -1330 -616 -1154
rect -674 -1342 -616 -1330
rect -416 -1154 -358 -1142
rect -416 -1330 -404 -1154
rect -370 -1330 -358 -1154
rect -416 -1342 -358 -1330
rect -158 -1154 -100 -1142
rect -158 -1330 -146 -1154
rect -112 -1330 -100 -1154
rect -158 -1342 -100 -1330
rect 100 -1154 158 -1142
rect 100 -1330 112 -1154
rect 146 -1330 158 -1154
rect 100 -1342 158 -1330
rect 358 -1154 416 -1142
rect 358 -1330 370 -1154
rect 404 -1330 416 -1154
rect 358 -1342 416 -1330
rect 616 -1154 674 -1142
rect 616 -1330 628 -1154
rect 662 -1330 674 -1154
rect 616 -1342 674 -1330
rect 874 -1154 932 -1142
rect 874 -1330 886 -1154
rect 920 -1330 932 -1154
rect 874 -1342 932 -1330
<< pdiffc >>
rect -920 1225 -886 1401
rect -662 1225 -628 1401
rect -404 1225 -370 1401
rect -146 1225 -112 1401
rect 112 1225 146 1401
rect 370 1225 404 1401
rect 628 1225 662 1401
rect 886 1225 920 1401
rect -920 860 -886 1036
rect -662 860 -628 1036
rect -404 860 -370 1036
rect -146 860 -112 1036
rect 112 860 146 1036
rect 370 860 404 1036
rect 628 860 662 1036
rect 886 860 920 1036
rect -920 495 -886 671
rect -662 495 -628 671
rect -404 495 -370 671
rect -146 495 -112 671
rect 112 495 146 671
rect 370 495 404 671
rect 628 495 662 671
rect 886 495 920 671
rect -920 130 -886 306
rect -662 130 -628 306
rect -404 130 -370 306
rect -146 130 -112 306
rect 112 130 146 306
rect 370 130 404 306
rect 628 130 662 306
rect 886 130 920 306
rect -920 -235 -886 -59
rect -662 -235 -628 -59
rect -404 -235 -370 -59
rect -146 -235 -112 -59
rect 112 -235 146 -59
rect 370 -235 404 -59
rect 628 -235 662 -59
rect 886 -235 920 -59
rect -920 -600 -886 -424
rect -662 -600 -628 -424
rect -404 -600 -370 -424
rect -146 -600 -112 -424
rect 112 -600 146 -424
rect 370 -600 404 -424
rect 628 -600 662 -424
rect 886 -600 920 -424
rect -920 -965 -886 -789
rect -662 -965 -628 -789
rect -404 -965 -370 -789
rect -146 -965 -112 -789
rect 112 -965 146 -789
rect 370 -965 404 -789
rect 628 -965 662 -789
rect 886 -965 920 -789
rect -920 -1330 -886 -1154
rect -662 -1330 -628 -1154
rect -404 -1330 -370 -1154
rect -146 -1330 -112 -1154
rect 112 -1330 146 -1154
rect 370 -1330 404 -1154
rect 628 -1330 662 -1154
rect 886 -1330 920 -1154
<< poly >>
rect -874 1413 -674 1439
rect -616 1413 -416 1439
rect -358 1413 -158 1439
rect -100 1413 100 1439
rect 158 1413 358 1439
rect 416 1413 616 1439
rect 674 1413 874 1439
rect -874 1166 -674 1213
rect -874 1132 -858 1166
rect -690 1132 -674 1166
rect -874 1116 -674 1132
rect -616 1166 -416 1213
rect -616 1132 -600 1166
rect -432 1132 -416 1166
rect -616 1116 -416 1132
rect -358 1166 -158 1213
rect -358 1132 -342 1166
rect -174 1132 -158 1166
rect -358 1116 -158 1132
rect -100 1166 100 1213
rect -100 1132 -84 1166
rect 84 1132 100 1166
rect -100 1116 100 1132
rect 158 1166 358 1213
rect 158 1132 174 1166
rect 342 1132 358 1166
rect 158 1116 358 1132
rect 416 1166 616 1213
rect 416 1132 432 1166
rect 600 1132 616 1166
rect 416 1116 616 1132
rect 674 1166 874 1213
rect 674 1132 690 1166
rect 858 1132 874 1166
rect 674 1116 874 1132
rect -874 1048 -674 1074
rect -616 1048 -416 1074
rect -358 1048 -158 1074
rect -100 1048 100 1074
rect 158 1048 358 1074
rect 416 1048 616 1074
rect 674 1048 874 1074
rect -874 801 -674 848
rect -874 767 -858 801
rect -690 767 -674 801
rect -874 751 -674 767
rect -616 801 -416 848
rect -616 767 -600 801
rect -432 767 -416 801
rect -616 751 -416 767
rect -358 801 -158 848
rect -358 767 -342 801
rect -174 767 -158 801
rect -358 751 -158 767
rect -100 801 100 848
rect -100 767 -84 801
rect 84 767 100 801
rect -100 751 100 767
rect 158 801 358 848
rect 158 767 174 801
rect 342 767 358 801
rect 158 751 358 767
rect 416 801 616 848
rect 416 767 432 801
rect 600 767 616 801
rect 416 751 616 767
rect 674 801 874 848
rect 674 767 690 801
rect 858 767 874 801
rect 674 751 874 767
rect -874 683 -674 709
rect -616 683 -416 709
rect -358 683 -158 709
rect -100 683 100 709
rect 158 683 358 709
rect 416 683 616 709
rect 674 683 874 709
rect -874 436 -674 483
rect -874 402 -858 436
rect -690 402 -674 436
rect -874 386 -674 402
rect -616 436 -416 483
rect -616 402 -600 436
rect -432 402 -416 436
rect -616 386 -416 402
rect -358 436 -158 483
rect -358 402 -342 436
rect -174 402 -158 436
rect -358 386 -158 402
rect -100 436 100 483
rect -100 402 -84 436
rect 84 402 100 436
rect -100 386 100 402
rect 158 436 358 483
rect 158 402 174 436
rect 342 402 358 436
rect 158 386 358 402
rect 416 436 616 483
rect 416 402 432 436
rect 600 402 616 436
rect 416 386 616 402
rect 674 436 874 483
rect 674 402 690 436
rect 858 402 874 436
rect 674 386 874 402
rect -874 318 -674 344
rect -616 318 -416 344
rect -358 318 -158 344
rect -100 318 100 344
rect 158 318 358 344
rect 416 318 616 344
rect 674 318 874 344
rect -874 71 -674 118
rect -874 37 -858 71
rect -690 37 -674 71
rect -874 21 -674 37
rect -616 71 -416 118
rect -616 37 -600 71
rect -432 37 -416 71
rect -616 21 -416 37
rect -358 71 -158 118
rect -358 37 -342 71
rect -174 37 -158 71
rect -358 21 -158 37
rect -100 71 100 118
rect -100 37 -84 71
rect 84 37 100 71
rect -100 21 100 37
rect 158 71 358 118
rect 158 37 174 71
rect 342 37 358 71
rect 158 21 358 37
rect 416 71 616 118
rect 416 37 432 71
rect 600 37 616 71
rect 416 21 616 37
rect 674 71 874 118
rect 674 37 690 71
rect 858 37 874 71
rect 674 21 874 37
rect -874 -47 -674 -21
rect -616 -47 -416 -21
rect -358 -47 -158 -21
rect -100 -47 100 -21
rect 158 -47 358 -21
rect 416 -47 616 -21
rect 674 -47 874 -21
rect -874 -294 -674 -247
rect -874 -328 -858 -294
rect -690 -328 -674 -294
rect -874 -344 -674 -328
rect -616 -294 -416 -247
rect -616 -328 -600 -294
rect -432 -328 -416 -294
rect -616 -344 -416 -328
rect -358 -294 -158 -247
rect -358 -328 -342 -294
rect -174 -328 -158 -294
rect -358 -344 -158 -328
rect -100 -294 100 -247
rect -100 -328 -84 -294
rect 84 -328 100 -294
rect -100 -344 100 -328
rect 158 -294 358 -247
rect 158 -328 174 -294
rect 342 -328 358 -294
rect 158 -344 358 -328
rect 416 -294 616 -247
rect 416 -328 432 -294
rect 600 -328 616 -294
rect 416 -344 616 -328
rect 674 -294 874 -247
rect 674 -328 690 -294
rect 858 -328 874 -294
rect 674 -344 874 -328
rect -874 -412 -674 -386
rect -616 -412 -416 -386
rect -358 -412 -158 -386
rect -100 -412 100 -386
rect 158 -412 358 -386
rect 416 -412 616 -386
rect 674 -412 874 -386
rect -874 -659 -674 -612
rect -874 -693 -858 -659
rect -690 -693 -674 -659
rect -874 -709 -674 -693
rect -616 -659 -416 -612
rect -616 -693 -600 -659
rect -432 -693 -416 -659
rect -616 -709 -416 -693
rect -358 -659 -158 -612
rect -358 -693 -342 -659
rect -174 -693 -158 -659
rect -358 -709 -158 -693
rect -100 -659 100 -612
rect -100 -693 -84 -659
rect 84 -693 100 -659
rect -100 -709 100 -693
rect 158 -659 358 -612
rect 158 -693 174 -659
rect 342 -693 358 -659
rect 158 -709 358 -693
rect 416 -659 616 -612
rect 416 -693 432 -659
rect 600 -693 616 -659
rect 416 -709 616 -693
rect 674 -659 874 -612
rect 674 -693 690 -659
rect 858 -693 874 -659
rect 674 -709 874 -693
rect -874 -777 -674 -751
rect -616 -777 -416 -751
rect -358 -777 -158 -751
rect -100 -777 100 -751
rect 158 -777 358 -751
rect 416 -777 616 -751
rect 674 -777 874 -751
rect -874 -1024 -674 -977
rect -874 -1058 -858 -1024
rect -690 -1058 -674 -1024
rect -874 -1074 -674 -1058
rect -616 -1024 -416 -977
rect -616 -1058 -600 -1024
rect -432 -1058 -416 -1024
rect -616 -1074 -416 -1058
rect -358 -1024 -158 -977
rect -358 -1058 -342 -1024
rect -174 -1058 -158 -1024
rect -358 -1074 -158 -1058
rect -100 -1024 100 -977
rect -100 -1058 -84 -1024
rect 84 -1058 100 -1024
rect -100 -1074 100 -1058
rect 158 -1024 358 -977
rect 158 -1058 174 -1024
rect 342 -1058 358 -1024
rect 158 -1074 358 -1058
rect 416 -1024 616 -977
rect 416 -1058 432 -1024
rect 600 -1058 616 -1024
rect 416 -1074 616 -1058
rect 674 -1024 874 -977
rect 674 -1058 690 -1024
rect 858 -1058 874 -1024
rect 674 -1074 874 -1058
rect -874 -1142 -674 -1116
rect -616 -1142 -416 -1116
rect -358 -1142 -158 -1116
rect -100 -1142 100 -1116
rect 158 -1142 358 -1116
rect 416 -1142 616 -1116
rect 674 -1142 874 -1116
rect -874 -1389 -674 -1342
rect -874 -1423 -858 -1389
rect -690 -1423 -674 -1389
rect -874 -1439 -674 -1423
rect -616 -1389 -416 -1342
rect -616 -1423 -600 -1389
rect -432 -1423 -416 -1389
rect -616 -1439 -416 -1423
rect -358 -1389 -158 -1342
rect -358 -1423 -342 -1389
rect -174 -1423 -158 -1389
rect -358 -1439 -158 -1423
rect -100 -1389 100 -1342
rect -100 -1423 -84 -1389
rect 84 -1423 100 -1389
rect -100 -1439 100 -1423
rect 158 -1389 358 -1342
rect 158 -1423 174 -1389
rect 342 -1423 358 -1389
rect 158 -1439 358 -1423
rect 416 -1389 616 -1342
rect 416 -1423 432 -1389
rect 600 -1423 616 -1389
rect 416 -1439 616 -1423
rect 674 -1389 874 -1342
rect 674 -1423 690 -1389
rect 858 -1423 874 -1389
rect 674 -1439 874 -1423
<< polycont >>
rect -858 1132 -690 1166
rect -600 1132 -432 1166
rect -342 1132 -174 1166
rect -84 1132 84 1166
rect 174 1132 342 1166
rect 432 1132 600 1166
rect 690 1132 858 1166
rect -858 767 -690 801
rect -600 767 -432 801
rect -342 767 -174 801
rect -84 767 84 801
rect 174 767 342 801
rect 432 767 600 801
rect 690 767 858 801
rect -858 402 -690 436
rect -600 402 -432 436
rect -342 402 -174 436
rect -84 402 84 436
rect 174 402 342 436
rect 432 402 600 436
rect 690 402 858 436
rect -858 37 -690 71
rect -600 37 -432 71
rect -342 37 -174 71
rect -84 37 84 71
rect 174 37 342 71
rect 432 37 600 71
rect 690 37 858 71
rect -858 -328 -690 -294
rect -600 -328 -432 -294
rect -342 -328 -174 -294
rect -84 -328 84 -294
rect 174 -328 342 -294
rect 432 -328 600 -294
rect 690 -328 858 -294
rect -858 -693 -690 -659
rect -600 -693 -432 -659
rect -342 -693 -174 -659
rect -84 -693 84 -659
rect 174 -693 342 -659
rect 432 -693 600 -659
rect 690 -693 858 -659
rect -858 -1058 -690 -1024
rect -600 -1058 -432 -1024
rect -342 -1058 -174 -1024
rect -84 -1058 84 -1024
rect 174 -1058 342 -1024
rect 432 -1058 600 -1024
rect 690 -1058 858 -1024
rect -858 -1423 -690 -1389
rect -600 -1423 -432 -1389
rect -342 -1423 -174 -1389
rect -84 -1423 84 -1389
rect 174 -1423 342 -1389
rect 432 -1423 600 -1389
rect 690 -1423 858 -1389
<< locali >>
rect -920 1401 -886 1417
rect -920 1209 -886 1225
rect -662 1401 -628 1417
rect -662 1209 -628 1225
rect -404 1401 -370 1417
rect -404 1209 -370 1225
rect -146 1401 -112 1417
rect -146 1209 -112 1225
rect 112 1401 146 1417
rect 112 1209 146 1225
rect 370 1401 404 1417
rect 370 1209 404 1225
rect 628 1401 662 1417
rect 628 1209 662 1225
rect 886 1401 920 1417
rect 886 1209 920 1225
rect -874 1132 -858 1166
rect -690 1132 -674 1166
rect -616 1132 -600 1166
rect -432 1132 -416 1166
rect -358 1132 -342 1166
rect -174 1132 -158 1166
rect -100 1132 -84 1166
rect 84 1132 100 1166
rect 158 1132 174 1166
rect 342 1132 358 1166
rect 416 1132 432 1166
rect 600 1132 616 1166
rect 674 1132 690 1166
rect 858 1132 874 1166
rect -920 1036 -886 1052
rect -920 844 -886 860
rect -662 1036 -628 1052
rect -662 844 -628 860
rect -404 1036 -370 1052
rect -404 844 -370 860
rect -146 1036 -112 1052
rect -146 844 -112 860
rect 112 1036 146 1052
rect 112 844 146 860
rect 370 1036 404 1052
rect 370 844 404 860
rect 628 1036 662 1052
rect 628 844 662 860
rect 886 1036 920 1052
rect 886 844 920 860
rect -874 767 -858 801
rect -690 767 -674 801
rect -616 767 -600 801
rect -432 767 -416 801
rect -358 767 -342 801
rect -174 767 -158 801
rect -100 767 -84 801
rect 84 767 100 801
rect 158 767 174 801
rect 342 767 358 801
rect 416 767 432 801
rect 600 767 616 801
rect 674 767 690 801
rect 858 767 874 801
rect -920 671 -886 687
rect -920 479 -886 495
rect -662 671 -628 687
rect -662 479 -628 495
rect -404 671 -370 687
rect -404 479 -370 495
rect -146 671 -112 687
rect -146 479 -112 495
rect 112 671 146 687
rect 112 479 146 495
rect 370 671 404 687
rect 370 479 404 495
rect 628 671 662 687
rect 628 479 662 495
rect 886 671 920 687
rect 886 479 920 495
rect -874 402 -858 436
rect -690 402 -674 436
rect -616 402 -600 436
rect -432 402 -416 436
rect -358 402 -342 436
rect -174 402 -158 436
rect -100 402 -84 436
rect 84 402 100 436
rect 158 402 174 436
rect 342 402 358 436
rect 416 402 432 436
rect 600 402 616 436
rect 674 402 690 436
rect 858 402 874 436
rect -920 306 -886 322
rect -920 114 -886 130
rect -662 306 -628 322
rect -662 114 -628 130
rect -404 306 -370 322
rect -404 114 -370 130
rect -146 306 -112 322
rect -146 114 -112 130
rect 112 306 146 322
rect 112 114 146 130
rect 370 306 404 322
rect 370 114 404 130
rect 628 306 662 322
rect 628 114 662 130
rect 886 306 920 322
rect 886 114 920 130
rect -874 37 -858 71
rect -690 37 -674 71
rect -616 37 -600 71
rect -432 37 -416 71
rect -358 37 -342 71
rect -174 37 -158 71
rect -100 37 -84 71
rect 84 37 100 71
rect 158 37 174 71
rect 342 37 358 71
rect 416 37 432 71
rect 600 37 616 71
rect 674 37 690 71
rect 858 37 874 71
rect -920 -59 -886 -43
rect -920 -251 -886 -235
rect -662 -59 -628 -43
rect -662 -251 -628 -235
rect -404 -59 -370 -43
rect -404 -251 -370 -235
rect -146 -59 -112 -43
rect -146 -251 -112 -235
rect 112 -59 146 -43
rect 112 -251 146 -235
rect 370 -59 404 -43
rect 370 -251 404 -235
rect 628 -59 662 -43
rect 628 -251 662 -235
rect 886 -59 920 -43
rect 886 -251 920 -235
rect -874 -328 -858 -294
rect -690 -328 -674 -294
rect -616 -328 -600 -294
rect -432 -328 -416 -294
rect -358 -328 -342 -294
rect -174 -328 -158 -294
rect -100 -328 -84 -294
rect 84 -328 100 -294
rect 158 -328 174 -294
rect 342 -328 358 -294
rect 416 -328 432 -294
rect 600 -328 616 -294
rect 674 -328 690 -294
rect 858 -328 874 -294
rect -920 -424 -886 -408
rect -920 -616 -886 -600
rect -662 -424 -628 -408
rect -662 -616 -628 -600
rect -404 -424 -370 -408
rect -404 -616 -370 -600
rect -146 -424 -112 -408
rect -146 -616 -112 -600
rect 112 -424 146 -408
rect 112 -616 146 -600
rect 370 -424 404 -408
rect 370 -616 404 -600
rect 628 -424 662 -408
rect 628 -616 662 -600
rect 886 -424 920 -408
rect 886 -616 920 -600
rect -874 -693 -858 -659
rect -690 -693 -674 -659
rect -616 -693 -600 -659
rect -432 -693 -416 -659
rect -358 -693 -342 -659
rect -174 -693 -158 -659
rect -100 -693 -84 -659
rect 84 -693 100 -659
rect 158 -693 174 -659
rect 342 -693 358 -659
rect 416 -693 432 -659
rect 600 -693 616 -659
rect 674 -693 690 -659
rect 858 -693 874 -659
rect -920 -789 -886 -773
rect -920 -981 -886 -965
rect -662 -789 -628 -773
rect -662 -981 -628 -965
rect -404 -789 -370 -773
rect -404 -981 -370 -965
rect -146 -789 -112 -773
rect -146 -981 -112 -965
rect 112 -789 146 -773
rect 112 -981 146 -965
rect 370 -789 404 -773
rect 370 -981 404 -965
rect 628 -789 662 -773
rect 628 -981 662 -965
rect 886 -789 920 -773
rect 886 -981 920 -965
rect -874 -1058 -858 -1024
rect -690 -1058 -674 -1024
rect -616 -1058 -600 -1024
rect -432 -1058 -416 -1024
rect -358 -1058 -342 -1024
rect -174 -1058 -158 -1024
rect -100 -1058 -84 -1024
rect 84 -1058 100 -1024
rect 158 -1058 174 -1024
rect 342 -1058 358 -1024
rect 416 -1058 432 -1024
rect 600 -1058 616 -1024
rect 674 -1058 690 -1024
rect 858 -1058 874 -1024
rect -920 -1154 -886 -1138
rect -920 -1346 -886 -1330
rect -662 -1154 -628 -1138
rect -662 -1346 -628 -1330
rect -404 -1154 -370 -1138
rect -404 -1346 -370 -1330
rect -146 -1154 -112 -1138
rect -146 -1346 -112 -1330
rect 112 -1154 146 -1138
rect 112 -1346 146 -1330
rect 370 -1154 404 -1138
rect 370 -1346 404 -1330
rect 628 -1154 662 -1138
rect 628 -1346 662 -1330
rect 886 -1154 920 -1138
rect 886 -1346 920 -1330
rect -874 -1423 -858 -1389
rect -690 -1423 -674 -1389
rect -616 -1423 -600 -1389
rect -432 -1423 -416 -1389
rect -358 -1423 -342 -1389
rect -174 -1423 -158 -1389
rect -100 -1423 -84 -1389
rect 84 -1423 100 -1389
rect 158 -1423 174 -1389
rect 342 -1423 358 -1389
rect 416 -1423 432 -1389
rect 600 -1423 616 -1389
rect 674 -1423 690 -1389
rect 858 -1423 874 -1389
<< viali >>
rect -920 1225 -886 1401
rect -662 1225 -628 1401
rect -404 1225 -370 1401
rect -146 1225 -112 1401
rect 112 1225 146 1401
rect 370 1225 404 1401
rect 628 1225 662 1401
rect 886 1225 920 1401
rect -858 1132 -690 1166
rect -600 1132 -432 1166
rect -342 1132 -174 1166
rect -84 1132 84 1166
rect 174 1132 342 1166
rect 432 1132 600 1166
rect 690 1132 858 1166
rect -920 860 -886 1036
rect -662 860 -628 1036
rect -404 860 -370 1036
rect -146 860 -112 1036
rect 112 860 146 1036
rect 370 860 404 1036
rect 628 860 662 1036
rect 886 860 920 1036
rect -858 767 -690 801
rect -600 767 -432 801
rect -342 767 -174 801
rect -84 767 84 801
rect 174 767 342 801
rect 432 767 600 801
rect 690 767 858 801
rect -920 495 -886 671
rect -662 495 -628 671
rect -404 495 -370 671
rect -146 495 -112 671
rect 112 495 146 671
rect 370 495 404 671
rect 628 495 662 671
rect 886 495 920 671
rect -858 402 -690 436
rect -600 402 -432 436
rect -342 402 -174 436
rect -84 402 84 436
rect 174 402 342 436
rect 432 402 600 436
rect 690 402 858 436
rect -920 130 -886 306
rect -662 130 -628 306
rect -404 130 -370 306
rect -146 130 -112 306
rect 112 130 146 306
rect 370 130 404 306
rect 628 130 662 306
rect 886 130 920 306
rect -858 37 -690 71
rect -600 37 -432 71
rect -342 37 -174 71
rect -84 37 84 71
rect 174 37 342 71
rect 432 37 600 71
rect 690 37 858 71
rect -920 -235 -886 -59
rect -662 -235 -628 -59
rect -404 -235 -370 -59
rect -146 -235 -112 -59
rect 112 -235 146 -59
rect 370 -235 404 -59
rect 628 -235 662 -59
rect 886 -235 920 -59
rect -858 -328 -690 -294
rect -600 -328 -432 -294
rect -342 -328 -174 -294
rect -84 -328 84 -294
rect 174 -328 342 -294
rect 432 -328 600 -294
rect 690 -328 858 -294
rect -920 -600 -886 -424
rect -662 -600 -628 -424
rect -404 -600 -370 -424
rect -146 -600 -112 -424
rect 112 -600 146 -424
rect 370 -600 404 -424
rect 628 -600 662 -424
rect 886 -600 920 -424
rect -858 -693 -690 -659
rect -600 -693 -432 -659
rect -342 -693 -174 -659
rect -84 -693 84 -659
rect 174 -693 342 -659
rect 432 -693 600 -659
rect 690 -693 858 -659
rect -920 -965 -886 -789
rect -662 -965 -628 -789
rect -404 -965 -370 -789
rect -146 -965 -112 -789
rect 112 -965 146 -789
rect 370 -965 404 -789
rect 628 -965 662 -789
rect 886 -965 920 -789
rect -858 -1058 -690 -1024
rect -600 -1058 -432 -1024
rect -342 -1058 -174 -1024
rect -84 -1058 84 -1024
rect 174 -1058 342 -1024
rect 432 -1058 600 -1024
rect 690 -1058 858 -1024
rect -920 -1330 -886 -1154
rect -662 -1330 -628 -1154
rect -404 -1330 -370 -1154
rect -146 -1330 -112 -1154
rect 112 -1330 146 -1154
rect 370 -1330 404 -1154
rect 628 -1330 662 -1154
rect 886 -1330 920 -1154
rect -858 -1423 -690 -1389
rect -600 -1423 -432 -1389
rect -342 -1423 -174 -1389
rect -84 -1423 84 -1389
rect 174 -1423 342 -1389
rect 432 -1423 600 -1389
rect 690 -1423 858 -1389
<< metal1 >>
rect -926 1401 -880 1413
rect -926 1225 -920 1401
rect -886 1225 -880 1401
rect -926 1213 -880 1225
rect -668 1401 -622 1413
rect -668 1225 -662 1401
rect -628 1225 -622 1401
rect -668 1213 -622 1225
rect -410 1401 -364 1413
rect -410 1225 -404 1401
rect -370 1225 -364 1401
rect -410 1213 -364 1225
rect -152 1401 -106 1413
rect -152 1225 -146 1401
rect -112 1225 -106 1401
rect -152 1213 -106 1225
rect 106 1401 152 1413
rect 106 1225 112 1401
rect 146 1225 152 1401
rect 106 1213 152 1225
rect 364 1401 410 1413
rect 364 1225 370 1401
rect 404 1225 410 1401
rect 364 1213 410 1225
rect 622 1401 668 1413
rect 622 1225 628 1401
rect 662 1225 668 1401
rect 622 1213 668 1225
rect 880 1401 926 1413
rect 880 1225 886 1401
rect 920 1225 926 1401
rect 880 1213 926 1225
rect -870 1166 -678 1172
rect -870 1132 -858 1166
rect -690 1132 -678 1166
rect -870 1126 -678 1132
rect -612 1166 -420 1172
rect -612 1132 -600 1166
rect -432 1132 -420 1166
rect -612 1126 -420 1132
rect -354 1166 -162 1172
rect -354 1132 -342 1166
rect -174 1132 -162 1166
rect -354 1126 -162 1132
rect -96 1166 96 1172
rect -96 1132 -84 1166
rect 84 1132 96 1166
rect -96 1126 96 1132
rect 162 1166 354 1172
rect 162 1132 174 1166
rect 342 1132 354 1166
rect 162 1126 354 1132
rect 420 1166 612 1172
rect 420 1132 432 1166
rect 600 1132 612 1166
rect 420 1126 612 1132
rect 678 1166 870 1172
rect 678 1132 690 1166
rect 858 1132 870 1166
rect 678 1126 870 1132
rect -926 1036 -880 1048
rect -926 860 -920 1036
rect -886 860 -880 1036
rect -926 848 -880 860
rect -668 1036 -622 1048
rect -668 860 -662 1036
rect -628 860 -622 1036
rect -668 848 -622 860
rect -410 1036 -364 1048
rect -410 860 -404 1036
rect -370 860 -364 1036
rect -410 848 -364 860
rect -152 1036 -106 1048
rect -152 860 -146 1036
rect -112 860 -106 1036
rect -152 848 -106 860
rect 106 1036 152 1048
rect 106 860 112 1036
rect 146 860 152 1036
rect 106 848 152 860
rect 364 1036 410 1048
rect 364 860 370 1036
rect 404 860 410 1036
rect 364 848 410 860
rect 622 1036 668 1048
rect 622 860 628 1036
rect 662 860 668 1036
rect 622 848 668 860
rect 880 1036 926 1048
rect 880 860 886 1036
rect 920 860 926 1036
rect 880 848 926 860
rect -870 801 -678 807
rect -870 767 -858 801
rect -690 767 -678 801
rect -870 761 -678 767
rect -612 801 -420 807
rect -612 767 -600 801
rect -432 767 -420 801
rect -612 761 -420 767
rect -354 801 -162 807
rect -354 767 -342 801
rect -174 767 -162 801
rect -354 761 -162 767
rect -96 801 96 807
rect -96 767 -84 801
rect 84 767 96 801
rect -96 761 96 767
rect 162 801 354 807
rect 162 767 174 801
rect 342 767 354 801
rect 162 761 354 767
rect 420 801 612 807
rect 420 767 432 801
rect 600 767 612 801
rect 420 761 612 767
rect 678 801 870 807
rect 678 767 690 801
rect 858 767 870 801
rect 678 761 870 767
rect -926 671 -880 683
rect -926 495 -920 671
rect -886 495 -880 671
rect -926 483 -880 495
rect -668 671 -622 683
rect -668 495 -662 671
rect -628 495 -622 671
rect -668 483 -622 495
rect -410 671 -364 683
rect -410 495 -404 671
rect -370 495 -364 671
rect -410 483 -364 495
rect -152 671 -106 683
rect -152 495 -146 671
rect -112 495 -106 671
rect -152 483 -106 495
rect 106 671 152 683
rect 106 495 112 671
rect 146 495 152 671
rect 106 483 152 495
rect 364 671 410 683
rect 364 495 370 671
rect 404 495 410 671
rect 364 483 410 495
rect 622 671 668 683
rect 622 495 628 671
rect 662 495 668 671
rect 622 483 668 495
rect 880 671 926 683
rect 880 495 886 671
rect 920 495 926 671
rect 880 483 926 495
rect -870 436 -678 442
rect -870 402 -858 436
rect -690 402 -678 436
rect -870 396 -678 402
rect -612 436 -420 442
rect -612 402 -600 436
rect -432 402 -420 436
rect -612 396 -420 402
rect -354 436 -162 442
rect -354 402 -342 436
rect -174 402 -162 436
rect -354 396 -162 402
rect -96 436 96 442
rect -96 402 -84 436
rect 84 402 96 436
rect -96 396 96 402
rect 162 436 354 442
rect 162 402 174 436
rect 342 402 354 436
rect 162 396 354 402
rect 420 436 612 442
rect 420 402 432 436
rect 600 402 612 436
rect 420 396 612 402
rect 678 436 870 442
rect 678 402 690 436
rect 858 402 870 436
rect 678 396 870 402
rect -926 306 -880 318
rect -926 130 -920 306
rect -886 130 -880 306
rect -926 118 -880 130
rect -668 306 -622 318
rect -668 130 -662 306
rect -628 130 -622 306
rect -668 118 -622 130
rect -410 306 -364 318
rect -410 130 -404 306
rect -370 130 -364 306
rect -410 118 -364 130
rect -152 306 -106 318
rect -152 130 -146 306
rect -112 130 -106 306
rect -152 118 -106 130
rect 106 306 152 318
rect 106 130 112 306
rect 146 130 152 306
rect 106 118 152 130
rect 364 306 410 318
rect 364 130 370 306
rect 404 130 410 306
rect 364 118 410 130
rect 622 306 668 318
rect 622 130 628 306
rect 662 130 668 306
rect 622 118 668 130
rect 880 306 926 318
rect 880 130 886 306
rect 920 130 926 306
rect 880 118 926 130
rect -870 71 -678 77
rect -870 37 -858 71
rect -690 37 -678 71
rect -870 31 -678 37
rect -612 71 -420 77
rect -612 37 -600 71
rect -432 37 -420 71
rect -612 31 -420 37
rect -354 71 -162 77
rect -354 37 -342 71
rect -174 37 -162 71
rect -354 31 -162 37
rect -96 71 96 77
rect -96 37 -84 71
rect 84 37 96 71
rect -96 31 96 37
rect 162 71 354 77
rect 162 37 174 71
rect 342 37 354 71
rect 162 31 354 37
rect 420 71 612 77
rect 420 37 432 71
rect 600 37 612 71
rect 420 31 612 37
rect 678 71 870 77
rect 678 37 690 71
rect 858 37 870 71
rect 678 31 870 37
rect -926 -59 -880 -47
rect -926 -235 -920 -59
rect -886 -235 -880 -59
rect -926 -247 -880 -235
rect -668 -59 -622 -47
rect -668 -235 -662 -59
rect -628 -235 -622 -59
rect -668 -247 -622 -235
rect -410 -59 -364 -47
rect -410 -235 -404 -59
rect -370 -235 -364 -59
rect -410 -247 -364 -235
rect -152 -59 -106 -47
rect -152 -235 -146 -59
rect -112 -235 -106 -59
rect -152 -247 -106 -235
rect 106 -59 152 -47
rect 106 -235 112 -59
rect 146 -235 152 -59
rect 106 -247 152 -235
rect 364 -59 410 -47
rect 364 -235 370 -59
rect 404 -235 410 -59
rect 364 -247 410 -235
rect 622 -59 668 -47
rect 622 -235 628 -59
rect 662 -235 668 -59
rect 622 -247 668 -235
rect 880 -59 926 -47
rect 880 -235 886 -59
rect 920 -235 926 -59
rect 880 -247 926 -235
rect -870 -294 -678 -288
rect -870 -328 -858 -294
rect -690 -328 -678 -294
rect -870 -334 -678 -328
rect -612 -294 -420 -288
rect -612 -328 -600 -294
rect -432 -328 -420 -294
rect -612 -334 -420 -328
rect -354 -294 -162 -288
rect -354 -328 -342 -294
rect -174 -328 -162 -294
rect -354 -334 -162 -328
rect -96 -294 96 -288
rect -96 -328 -84 -294
rect 84 -328 96 -294
rect -96 -334 96 -328
rect 162 -294 354 -288
rect 162 -328 174 -294
rect 342 -328 354 -294
rect 162 -334 354 -328
rect 420 -294 612 -288
rect 420 -328 432 -294
rect 600 -328 612 -294
rect 420 -334 612 -328
rect 678 -294 870 -288
rect 678 -328 690 -294
rect 858 -328 870 -294
rect 678 -334 870 -328
rect -926 -424 -880 -412
rect -926 -600 -920 -424
rect -886 -600 -880 -424
rect -926 -612 -880 -600
rect -668 -424 -622 -412
rect -668 -600 -662 -424
rect -628 -600 -622 -424
rect -668 -612 -622 -600
rect -410 -424 -364 -412
rect -410 -600 -404 -424
rect -370 -600 -364 -424
rect -410 -612 -364 -600
rect -152 -424 -106 -412
rect -152 -600 -146 -424
rect -112 -600 -106 -424
rect -152 -612 -106 -600
rect 106 -424 152 -412
rect 106 -600 112 -424
rect 146 -600 152 -424
rect 106 -612 152 -600
rect 364 -424 410 -412
rect 364 -600 370 -424
rect 404 -600 410 -424
rect 364 -612 410 -600
rect 622 -424 668 -412
rect 622 -600 628 -424
rect 662 -600 668 -424
rect 622 -612 668 -600
rect 880 -424 926 -412
rect 880 -600 886 -424
rect 920 -600 926 -424
rect 880 -612 926 -600
rect -870 -659 -678 -653
rect -870 -693 -858 -659
rect -690 -693 -678 -659
rect -870 -699 -678 -693
rect -612 -659 -420 -653
rect -612 -693 -600 -659
rect -432 -693 -420 -659
rect -612 -699 -420 -693
rect -354 -659 -162 -653
rect -354 -693 -342 -659
rect -174 -693 -162 -659
rect -354 -699 -162 -693
rect -96 -659 96 -653
rect -96 -693 -84 -659
rect 84 -693 96 -659
rect -96 -699 96 -693
rect 162 -659 354 -653
rect 162 -693 174 -659
rect 342 -693 354 -659
rect 162 -699 354 -693
rect 420 -659 612 -653
rect 420 -693 432 -659
rect 600 -693 612 -659
rect 420 -699 612 -693
rect 678 -659 870 -653
rect 678 -693 690 -659
rect 858 -693 870 -659
rect 678 -699 870 -693
rect -926 -789 -880 -777
rect -926 -965 -920 -789
rect -886 -965 -880 -789
rect -926 -977 -880 -965
rect -668 -789 -622 -777
rect -668 -965 -662 -789
rect -628 -965 -622 -789
rect -668 -977 -622 -965
rect -410 -789 -364 -777
rect -410 -965 -404 -789
rect -370 -965 -364 -789
rect -410 -977 -364 -965
rect -152 -789 -106 -777
rect -152 -965 -146 -789
rect -112 -965 -106 -789
rect -152 -977 -106 -965
rect 106 -789 152 -777
rect 106 -965 112 -789
rect 146 -965 152 -789
rect 106 -977 152 -965
rect 364 -789 410 -777
rect 364 -965 370 -789
rect 404 -965 410 -789
rect 364 -977 410 -965
rect 622 -789 668 -777
rect 622 -965 628 -789
rect 662 -965 668 -789
rect 622 -977 668 -965
rect 880 -789 926 -777
rect 880 -965 886 -789
rect 920 -965 926 -789
rect 880 -977 926 -965
rect -870 -1024 -678 -1018
rect -870 -1058 -858 -1024
rect -690 -1058 -678 -1024
rect -870 -1064 -678 -1058
rect -612 -1024 -420 -1018
rect -612 -1058 -600 -1024
rect -432 -1058 -420 -1024
rect -612 -1064 -420 -1058
rect -354 -1024 -162 -1018
rect -354 -1058 -342 -1024
rect -174 -1058 -162 -1024
rect -354 -1064 -162 -1058
rect -96 -1024 96 -1018
rect -96 -1058 -84 -1024
rect 84 -1058 96 -1024
rect -96 -1064 96 -1058
rect 162 -1024 354 -1018
rect 162 -1058 174 -1024
rect 342 -1058 354 -1024
rect 162 -1064 354 -1058
rect 420 -1024 612 -1018
rect 420 -1058 432 -1024
rect 600 -1058 612 -1024
rect 420 -1064 612 -1058
rect 678 -1024 870 -1018
rect 678 -1058 690 -1024
rect 858 -1058 870 -1024
rect 678 -1064 870 -1058
rect -926 -1154 -880 -1142
rect -926 -1330 -920 -1154
rect -886 -1330 -880 -1154
rect -926 -1342 -880 -1330
rect -668 -1154 -622 -1142
rect -668 -1330 -662 -1154
rect -628 -1330 -622 -1154
rect -668 -1342 -622 -1330
rect -410 -1154 -364 -1142
rect -410 -1330 -404 -1154
rect -370 -1330 -364 -1154
rect -410 -1342 -364 -1330
rect -152 -1154 -106 -1142
rect -152 -1330 -146 -1154
rect -112 -1330 -106 -1154
rect -152 -1342 -106 -1330
rect 106 -1154 152 -1142
rect 106 -1330 112 -1154
rect 146 -1330 152 -1154
rect 106 -1342 152 -1330
rect 364 -1154 410 -1142
rect 364 -1330 370 -1154
rect 404 -1330 410 -1154
rect 364 -1342 410 -1330
rect 622 -1154 668 -1142
rect 622 -1330 628 -1154
rect 662 -1330 668 -1154
rect 622 -1342 668 -1330
rect 880 -1154 926 -1142
rect 880 -1330 886 -1154
rect 920 -1330 926 -1154
rect 880 -1342 926 -1330
rect -870 -1389 -678 -1383
rect -870 -1423 -858 -1389
rect -690 -1423 -678 -1389
rect -870 -1429 -678 -1423
rect -612 -1389 -420 -1383
rect -612 -1423 -600 -1389
rect -432 -1423 -420 -1389
rect -612 -1429 -420 -1423
rect -354 -1389 -162 -1383
rect -354 -1423 -342 -1389
rect -174 -1423 -162 -1389
rect -354 -1429 -162 -1423
rect -96 -1389 96 -1383
rect -96 -1423 -84 -1389
rect 84 -1423 96 -1389
rect -96 -1429 96 -1423
rect 162 -1389 354 -1383
rect 162 -1423 174 -1389
rect 342 -1423 354 -1389
rect 162 -1429 354 -1423
rect 420 -1389 612 -1383
rect 420 -1423 432 -1389
rect 600 -1423 612 -1389
rect 420 -1429 612 -1423
rect 678 -1389 870 -1383
rect 678 -1423 690 -1389
rect 858 -1423 870 -1389
rect 678 -1429 870 -1423
<< properties >>
string gencell sky130_fd_pr__pfet_01v8_lvt
string library sky130
string parameters w 1 l 1 m 8 nf 7 diffcov 100 polycov 100 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 0 botc 1 poverlap 0 doverlap 1 lmin 0.35 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 0 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
