magic
tech sky130A
magscale 1 2
timestamp 1662665761
<< locali >>
rect 12290 11270 12670 11305
rect 12290 8660 12670 8695
rect 10175 7140 10215 8395
rect 11345 7140 11385 8395
rect 13575 7140 13615 8395
rect 14750 7140 14790 8395
rect 12290 6840 12670 6875
rect 12290 4230 12670 4265
<< metal2 >>
rect 12280 12036 14415 12111
rect 15735 12035 16085 12110
rect 15910 11825 15990 11835
rect 15910 11765 15920 11825
rect 15980 11765 15990 11825
rect 15910 11750 15990 11765
rect 15810 11460 15890 11470
rect 15810 11400 15820 11460
rect 15880 11400 15890 11460
rect 15810 11390 15890 11400
rect 9185 8265 10505 8275
rect 9185 8185 10425 8265
rect 10495 8185 10505 8265
rect 9185 8175 10505 8185
rect 10575 8145 10675 8330
rect 11130 8275 11230 8325
rect 13625 8320 13630 8380
rect 13625 8315 13635 8320
rect 14660 8370 14740 8395
rect 13695 8315 13705 8320
rect 13625 8305 13705 8315
rect 14660 8310 14670 8370
rect 14730 8310 14740 8370
rect 14660 8305 14740 8310
rect 10765 8265 15760 8275
rect 10765 8185 10775 8265
rect 10845 8185 12780 8265
rect 12860 8185 15760 8265
rect 10765 8175 15760 8185
rect 9185 8140 15760 8145
rect 9185 8055 14850 8140
rect 14930 8055 15760 8140
rect 9185 8045 15760 8055
rect 9185 8005 15760 8015
rect 9185 7925 10235 8005
rect 10295 7925 15760 8005
rect 9185 7915 15760 7925
rect 9185 7875 15760 7885
rect 9185 7795 11270 7875
rect 11330 7795 15760 7875
rect 9185 7785 15760 7795
rect 9185 7745 15760 7755
rect 9185 7665 13635 7745
rect 13695 7665 15760 7745
rect 9185 7655 15760 7665
rect 9185 7615 15760 7625
rect 9185 7535 14670 7615
rect 14730 7535 15760 7615
rect 9185 7525 15760 7535
rect 9180 7485 15760 7495
rect 9180 7405 12100 7485
rect 12190 7405 15760 7485
rect 9180 7395 15760 7405
rect 9175 7355 14190 7365
rect 9175 7275 9845 7355
rect 9925 7275 14120 7355
rect 14180 7275 14190 7355
rect 9175 7265 14190 7275
rect 10225 7225 10305 7235
rect 10225 7165 10235 7225
rect 10295 7165 10305 7225
rect 10225 7140 10305 7165
rect 11260 7225 11340 7235
rect 11260 7165 11270 7225
rect 11330 7165 11340 7225
rect 13755 7210 13830 7265
rect 14285 7215 14360 7395
rect 14460 7355 15760 7365
rect 14460 7275 14470 7355
rect 14530 7275 15760 7355
rect 14460 7265 15760 7275
rect 11260 7155 11340 7165
rect 15825 4175 15890 11390
rect 15815 4115 15825 4145
rect 15885 4115 15890 4175
rect 15815 4105 15890 4115
rect 15925 3770 15990 11750
rect 15910 3760 15990 3770
rect 15910 3700 15920 3760
rect 15980 3700 15990 3760
rect 15910 3685 15990 3700
rect 16020 3500 16085 12035
rect 12350 3425 13635 3500
rect 15730 3425 16085 3500
<< via2 >>
rect 15920 11765 15980 11825
rect 15820 11400 15880 11460
rect 10425 8185 10495 8265
rect 13635 8315 13695 8375
rect 14670 8310 14730 8370
rect 10775 8185 10845 8265
rect 12780 8185 12860 8265
rect 14850 8055 14930 8140
rect 10235 7925 10295 8005
rect 11270 7795 11330 7875
rect 13635 7665 13695 7745
rect 14670 7535 14730 7615
rect 12100 7405 12190 7485
rect 9845 7275 9925 7355
rect 14120 7275 14180 7355
rect 10235 7165 10295 7225
rect 11270 7165 11330 7225
rect 14470 7275 14530 7355
rect 15825 4115 15885 4175
rect 15920 3700 15980 3760
<< metal3 >>
rect 12355 11705 12775 12005
rect 15735 11825 15990 11835
rect 15735 11775 15920 11825
rect 15910 11765 15920 11775
rect 15980 11765 15990 11825
rect 15910 11750 15990 11765
rect 12350 11295 13540 11595
rect 15710 11460 15890 11470
rect 15710 11400 15820 11460
rect 15880 11400 15890 11460
rect 15710 11390 15890 11400
rect 10225 8005 10305 8460
rect 10415 8265 10855 8275
rect 10415 8185 10425 8265
rect 10495 8185 10775 8265
rect 10845 8185 10855 8265
rect 10415 8175 10855 8185
rect 10225 7925 10235 8005
rect 10295 7925 10305 8005
rect 9835 7355 9935 7365
rect 9835 7275 9845 7355
rect 9925 7275 9935 7355
rect 9835 6790 9935 7275
rect 10225 7225 10305 7925
rect 10225 7165 10235 7225
rect 10295 7165 10305 7225
rect 10225 7155 10305 7165
rect 11260 7875 11340 8445
rect 12770 8265 12870 8780
rect 12770 8185 12780 8265
rect 12860 8185 12870 8265
rect 12770 8175 12870 8185
rect 13625 8375 13705 8380
rect 13625 8315 13635 8375
rect 13695 8315 13705 8375
rect 11260 7795 11270 7875
rect 11330 7795 11340 7875
rect 11260 7225 11340 7795
rect 13625 7745 13705 8315
rect 13625 7665 13635 7745
rect 13695 7665 13705 7745
rect 11260 7165 11270 7225
rect 11330 7165 11340 7225
rect 11260 7155 11340 7165
rect 12095 7485 12195 7495
rect 12095 7405 12100 7485
rect 12190 7405 12195 7485
rect 12095 6790 12195 7405
rect 13625 7065 13705 7665
rect 14660 8370 14740 8380
rect 14660 8310 14670 8370
rect 14730 8310 14740 8370
rect 14660 7615 14740 8310
rect 14840 8140 14940 8740
rect 14840 8055 14850 8140
rect 14930 8055 14940 8140
rect 14840 8045 14940 8055
rect 14660 7535 14670 7615
rect 14730 7535 14740 7615
rect 14110 7355 14540 7365
rect 14110 7275 14120 7355
rect 14180 7275 14470 7355
rect 14530 7275 14540 7355
rect 14110 7265 14540 7275
rect 14660 7085 14740 7535
rect 12355 4075 13525 4240
rect 15725 4175 15890 4180
rect 15725 4120 15825 4175
rect 15750 4115 15825 4120
rect 15885 4115 15890 4175
rect 15750 4105 15890 4115
rect 12355 3940 13525 4005
rect 12355 3810 13525 3830
rect 12355 3550 12787 3810
rect 13317 3550 13525 3810
rect 15910 3760 15990 3770
rect 15910 3755 15920 3760
rect 15695 3700 15920 3755
rect 15980 3700 15990 3760
rect 15695 3685 15990 3700
rect 12355 3530 13525 3550
use core_osc_amp  X1
timestamp 1662515374
transform -1 0 14762 0 -1 12340
box 2396 230 5562 4020
use core_osc_amp  X2
timestamp 1662515374
transform -1 0 14762 0 1 3195
box 2396 230 5562 4020
use core_osc_amp  X3
timestamp 1662515374
transform -1 0 18162 0 1 3195
box 2396 230 5562 4020
use core_osc_amp  X4
timestamp 1662515374
transform -1 0 18162 0 -1 12340
box 2396 230 5562 4020
<< labels >>
rlabel metal2 9185 8045 14850 8145 1 S4A
rlabel metal2 9185 7915 10235 8015 1 S1B
rlabel metal2 9185 7785 11270 7885 1 S1A
rlabel metal2 9185 7655 13635 7755 1 S3B
rlabel metal2 9185 7525 14670 7625 1 S3A
rlabel metal2 9180 7395 12100 7495 1 S2A
rlabel metal2 9175 7265 9845 7365 1 S2B
rlabel metal2 14930 8045 15760 8145 1 S4A
rlabel metal2 10295 7915 15760 8015 1 S1B
rlabel metal2 11330 7785 15760 7885 1 S1A
rlabel metal2 13695 7655 15760 7755 1 S3B
rlabel metal2 14730 7525 15760 7625 1 S3A
rlabel metal2 12190 7395 15760 7495 1 S2A
rlabel metal2 14530 7265 15760 7365 1 S2B
rlabel metal2 9185 8175 10425 8275 1 S4B
rlabel metal2 12860 8175 15760 8275 1 S4B
rlabel metal2 16020 3425 16085 12110 1 BIAS
rlabel metal2 15925 3760 15990 11765 1 VDD
rlabel metal2 15825 4175 15890 11400 1 GND
rlabel locali 12290 8660 12670 8695 1 SUB
<< end >>
