magic
tech sky130A
magscale 1 2
timestamp 1662759368
<< pwell >>
rect -3223 -10998 3223 10998
<< psubdiff >>
rect -3187 10928 -3091 10962
rect 3091 10928 3187 10962
rect -3187 10866 -3153 10928
rect 3153 10866 3187 10928
rect -3187 -10928 -3153 -10866
rect 3153 -10928 3187 -10866
rect -3187 -10962 -3091 -10928
rect 3091 -10962 3187 -10928
<< psubdiffcont >>
rect -3091 10928 3091 10962
rect -3187 -10866 -3153 10866
rect 3153 -10866 3187 10866
rect -3091 -10962 3091 -10928
<< xpolycontact >>
rect -3057 10400 -1911 10832
rect -3057 -10832 -1911 -10400
rect -1815 10400 -669 10832
rect -1815 -10832 -669 -10400
rect -573 10400 573 10832
rect -573 -10832 573 -10400
rect 669 10400 1815 10832
rect 669 -10832 1815 -10400
rect 1911 10400 3057 10832
rect 1911 -10832 3057 -10400
<< xpolyres >>
rect -3057 -10400 -1911 10400
rect -1815 -10400 -669 10400
rect -573 -10400 573 10400
rect 669 -10400 1815 10400
rect 1911 -10400 3057 10400
<< locali >>
rect -3187 10928 -3091 10962
rect 3091 10928 3187 10962
rect -3187 10866 -3153 10928
rect 3153 10866 3187 10928
rect -3187 -10928 -3153 -10866
rect 3153 -10928 3187 -10866
rect -3187 -10962 -3091 -10928
rect 3091 -10962 3187 -10928
<< viali >>
rect -3041 10417 -1927 10814
rect -1799 10417 -685 10814
rect -557 10417 557 10814
rect 685 10417 1799 10814
rect 1927 10417 3041 10814
rect -3041 -10814 -1927 -10417
rect -1799 -10814 -685 -10417
rect -557 -10814 557 -10417
rect 685 -10814 1799 -10417
rect 1927 -10814 3041 -10417
<< metal1 >>
rect -3053 10814 -1915 10820
rect -3053 10417 -3041 10814
rect -1927 10417 -1915 10814
rect -3053 10411 -1915 10417
rect -1811 10814 -673 10820
rect -1811 10417 -1799 10814
rect -685 10417 -673 10814
rect -1811 10411 -673 10417
rect -569 10814 569 10820
rect -569 10417 -557 10814
rect 557 10417 569 10814
rect -569 10411 569 10417
rect 673 10814 1811 10820
rect 673 10417 685 10814
rect 1799 10417 1811 10814
rect 673 10411 1811 10417
rect 1915 10814 3053 10820
rect 1915 10417 1927 10814
rect 3041 10417 3053 10814
rect 1915 10411 3053 10417
rect -3053 -10417 -1915 -10411
rect -3053 -10814 -3041 -10417
rect -1927 -10814 -1915 -10417
rect -3053 -10820 -1915 -10814
rect -1811 -10417 -673 -10411
rect -1811 -10814 -1799 -10417
rect -685 -10814 -673 -10417
rect -1811 -10820 -673 -10814
rect -569 -10417 569 -10411
rect -569 -10814 -557 -10417
rect 557 -10814 569 -10417
rect -569 -10820 569 -10814
rect 673 -10417 1811 -10411
rect 673 -10814 685 -10417
rect 1799 -10814 1811 -10417
rect 673 -10820 1811 -10814
rect 1915 -10417 3053 -10411
rect 1915 -10814 1927 -10417
rect 3041 -10814 3053 -10417
rect 1915 -10820 3053 -10814
<< res5p73 >>
rect -3059 -10402 -1909 10402
rect -1817 -10402 -667 10402
rect -575 -10402 575 10402
rect 667 -10402 1817 10402
rect 1909 -10402 3059 10402
<< properties >>
string FIXED_BBOX -3170 -10945 3170 10945
string gencell sky130_fd_pr__res_xhigh_po_5p73
string library sky130
string parameters w 5.730 l 104 m 1 nx 5 wmin 5.730 lmin 0.50 rho 2000 val 36.365k dummy 0 dw 0.0 term 188.2 sterm 0.0 caplen 0 wmax 5.730 guard 1 glc 1 grc 1 gtc 1 gbc 1 compatible {sky130_fd_pr__res_xhigh_po_0p35  sky130_fd_pr__res_xhigh_po_0p69 sky130_fd_pr__res_xhigh_po_1p41  sky130_fd_pr__res_xhigh_po_2p85 sky130_fd_pr__res_xhigh_po_5p73} snake 0 full_metal 1 n_guard 0 hv_guard 0 vias 1 viagb 0 viagt 0 viagl 0 viagr 0
<< end >>
