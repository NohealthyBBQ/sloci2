magic
tech sky130A
magscale 1 2
timestamp 1662916051
<< pwell >>
rect -596 -679 596 679
<< nmoslvt >>
rect -400 -469 400 531
<< ndiff >>
rect -458 519 -400 531
rect -458 -457 -446 519
rect -412 -457 -400 519
rect -458 -469 -400 -457
rect 400 519 458 531
rect 400 -457 412 519
rect 446 -457 458 519
rect 400 -469 458 -457
<< ndiffc >>
rect -446 -457 -412 519
rect 412 -457 446 519
<< psubdiff >>
rect -560 609 560 643
rect -560 -609 -526 609
rect 526 -609 560 609
rect -560 -643 560 -609
<< poly >>
rect -400 531 400 557
rect -400 -507 400 -469
rect -400 -541 -384 -507
rect 384 -541 400 -507
rect -400 -557 400 -541
<< polycont >>
rect -384 -541 384 -507
<< locali >>
rect -560 609 560 643
rect -560 -609 -526 609
rect -446 519 -412 535
rect -446 -473 -412 -457
rect 412 519 446 535
rect 412 -473 446 -457
rect -400 -541 -384 -507
rect 384 -541 400 -507
rect 526 -609 560 609
rect -560 -643 560 -609
<< viali >>
rect -446 -457 -412 519
rect 412 -457 446 519
rect -384 -541 384 -507
<< metal1 >>
rect -452 519 -406 531
rect -452 -457 -446 519
rect -412 -457 -406 519
rect -452 -469 -406 -457
rect 406 519 452 531
rect 406 -457 412 519
rect 446 -457 452 519
rect 406 -469 452 -457
rect -396 -507 396 -501
rect -396 -541 -384 -507
rect 384 -541 396 -507
rect -396 -547 396 -541
<< properties >>
string FIXED_BBOX -543 -626 543 626
string gencell sky130_fd_pr__nfet_01v8_lvt
string library sky130
string parameters w 5 l 4 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 0 grc 0 gtc 0 gbc 0 tbcov 100 rlcov 100 topc 0 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
