magic
tech sky130A
magscale 1 2
timestamp 1672279567
<< error_p >>
rect -70 50 -10 6250
rect 10 50 70 6250
rect -70 -6250 -10 -50
rect 10 -6250 70 -50
<< metal3 >>
rect -6309 6222 -10 6250
rect -6309 78 -94 6222
rect -30 78 -10 6222
rect -6309 50 -10 78
rect 10 6222 6309 6250
rect 10 78 6225 6222
rect 6289 78 6309 6222
rect 10 50 6309 78
rect -6309 -78 -10 -50
rect -6309 -6222 -94 -78
rect -30 -6222 -10 -78
rect -6309 -6250 -10 -6222
rect 10 -78 6309 -50
rect 10 -6222 6225 -78
rect 6289 -6222 6309 -78
rect 10 -6250 6309 -6222
<< via3 >>
rect -94 78 -30 6222
rect 6225 78 6289 6222
rect -94 -6222 -30 -78
rect 6225 -6222 6289 -78
<< mimcap >>
rect -6209 6110 -209 6150
rect -6209 190 -6169 6110
rect -249 190 -209 6110
rect -6209 150 -209 190
rect 110 6110 6110 6150
rect 110 190 150 6110
rect 6070 190 6110 6110
rect 110 150 6110 190
rect -6209 -190 -209 -150
rect -6209 -6110 -6169 -190
rect -249 -6110 -209 -190
rect -6209 -6150 -209 -6110
rect 110 -190 6110 -150
rect 110 -6110 150 -190
rect 6070 -6110 6110 -190
rect 110 -6150 6110 -6110
<< mimcapcontact >>
rect -6169 190 -249 6110
rect 150 190 6070 6110
rect -6169 -6110 -249 -190
rect 150 -6110 6070 -190
<< metal4 >>
rect -3261 6111 -3157 6300
rect -141 6238 -37 6300
rect -141 6222 -14 6238
rect -6170 6110 -248 6111
rect -6170 190 -6169 6110
rect -249 190 -248 6110
rect -6170 189 -248 190
rect -3261 -189 -3157 189
rect -141 78 -94 6222
rect -30 78 -14 6222
rect 3058 6111 3162 6300
rect 6178 6238 6282 6300
rect 6178 6222 6305 6238
rect 149 6110 6071 6111
rect 149 190 150 6110
rect 6070 190 6071 6110
rect 149 189 6071 190
rect -141 62 -14 78
rect -141 -62 -37 62
rect -141 -78 -14 -62
rect -6170 -190 -248 -189
rect -6170 -6110 -6169 -190
rect -249 -6110 -248 -190
rect -6170 -6111 -248 -6110
rect -3261 -6300 -3157 -6111
rect -141 -6222 -94 -78
rect -30 -6222 -14 -78
rect 3058 -189 3162 189
rect 6178 78 6225 6222
rect 6289 78 6305 6222
rect 6178 62 6305 78
rect 6178 -62 6282 62
rect 6178 -78 6305 -62
rect 149 -190 6071 -189
rect 149 -6110 150 -190
rect 6070 -6110 6071 -190
rect 149 -6111 6071 -6110
rect -141 -6238 -14 -6222
rect -141 -6300 -37 -6238
rect 3058 -6300 3162 -6111
rect 6178 -6222 6225 -78
rect 6289 -6222 6305 -78
rect 6178 -6238 6305 -6222
rect 6178 -6300 6282 -6238
<< properties >>
string FIXED_BBOX 10 50 6210 6250
string gencell sky130_fd_pr__cap_mim_m3_1
string library sky130
string parameters w 30.0 l 30.0 val 1.822k carea 2.00 cperi 0.19 nx 2 ny 2 dummy 0 square 0 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 1 tconnect 1 ccov 100
<< end >>
