magic
tech sky130A
magscale 1 2
timestamp 1672438525
<< locali >>
rect 11660 5680 16200 5740
rect 11660 5420 16200 5490
rect 11660 5240 16210 5290
rect 11660 4990 16210 5040
rect 11720 4500 13100 4660
rect 14760 4500 16140 4660
rect 11720 4220 13100 4380
rect 14760 4220 16140 4380
rect 11660 3840 16210 3890
rect 11660 3590 16210 3640
rect 11670 3390 16220 3440
rect 11660 3140 16210 3190
<< metal1 >>
rect 17190 5680 17200 5980
rect 17560 5680 17570 5980
rect 13900 4010 13970 4560
rect 13890 3940 13900 4010
rect 13970 3940 13980 4010
rect 11790 2650 13030 2710
rect 12390 2560 12440 2650
rect 12370 2420 12380 2560
rect 12460 2420 12470 2560
rect 12390 2340 12440 2420
rect 11790 2290 13030 2340
rect 16620 -100 17600 -60
rect 16620 -360 16640 -100
rect 16960 -360 17600 -100
rect 38410 -320 38420 -100
rect 38800 -320 38810 -100
rect 16620 -380 17600 -360
rect 27630 -840 27640 -620
rect 28000 -840 28010 -620
<< via1 >>
rect 17200 5680 17560 5980
rect 13900 3940 13970 4010
rect 12380 2420 12460 2560
rect 16640 -360 16960 -100
rect 38420 -320 38800 -100
rect 27640 -840 28000 -620
<< metal2 >>
rect 17700 19880 18000 19900
rect 17700 19620 17720 19880
rect 17980 19620 18000 19880
rect 17700 19600 18000 19620
rect 16660 5980 17580 6000
rect 16660 5680 17200 5980
rect 17560 5680 17580 5980
rect 16660 5660 17580 5680
rect 16660 4580 17000 5660
rect 13100 4500 13600 4520
rect 13100 4380 13120 4500
rect 13240 4380 13600 4500
rect 13100 4360 13600 4380
rect 14000 4500 14200 4510
rect 14000 4290 14200 4300
rect 16660 4220 16680 4580
rect 16980 4220 17000 4580
rect 16660 4200 17000 4220
rect 11540 4010 13980 4020
rect 11540 3940 13900 4010
rect 13970 3940 13980 4010
rect 11540 3200 11620 3940
rect 13900 3930 13970 3940
rect 7300 3000 11620 3200
rect 11540 2540 11620 3000
rect 12380 2560 12460 2570
rect 11540 2420 12380 2540
rect 12380 2410 12460 2420
rect 1700 1860 1800 1870
rect 1700 1750 1800 1760
rect 2160 1860 2280 1880
rect 2160 1760 2170 1860
rect 2260 1760 2280 1860
rect 2160 20 2280 1760
rect 2160 -120 2180 20
rect 2260 -120 2280 20
rect 2160 -140 2280 -120
rect 16640 -100 16960 -90
rect 16640 -370 16960 -360
rect 38400 -100 38820 -80
rect 38400 -320 38420 -100
rect 38800 -320 38820 -100
rect 38400 -500 38820 -320
rect 27640 -620 38820 -500
rect 28000 -840 38820 -620
rect 27640 -960 38820 -840
<< via2 >>
rect 17720 19620 17980 19880
rect 13120 4380 13240 4500
rect 14000 4300 14200 4500
rect 16680 4220 16980 4580
rect 1700 1760 1800 1860
rect 2170 1760 2260 1860
rect 2180 -120 2260 20
rect 16640 -360 16960 -100
<< metal3 >>
rect 13000 19880 18000 19900
rect 13000 19620 17720 19880
rect 17980 19620 18000 19880
rect 13000 19600 18000 19620
rect 13000 6400 13400 19600
rect 13100 4500 13260 6400
rect 13100 4380 13120 4500
rect 13240 4380 13260 4500
rect 13100 4360 13260 4380
rect 13900 4580 17000 4600
rect 13900 4500 16680 4580
rect 13900 4300 14000 4500
rect 14200 4300 16680 4500
rect 13900 4220 16680 4300
rect 16980 4220 17000 4580
rect 13900 4200 17000 4220
rect 1690 1860 2270 1870
rect 1690 1760 1700 1860
rect 1800 1760 2170 1860
rect 2260 1760 2270 1860
rect 1690 1750 2270 1760
rect 16600 40 17000 4200
rect 2160 20 17000 40
rect 2160 -120 2180 20
rect 2260 -100 17000 20
rect 2260 -120 16640 -100
rect 2160 -140 16640 -120
rect 16600 -360 16640 -140
rect 16960 -360 17000 -100
rect 16600 -400 17000 -360
use XM_Rref  XM_Rref_0
timestamp 1662826901
transform 0 1 18173 1 0 1417
box -1417 -1173 5029 21223
use XM_current_gate_with_dummy  XM_current_gate_with_dummy_0
timestamp 1662842659
transform 1 0 11600 0 1 3924
box 0 -924 4660 1954
use XM_output_mirr_combined_with_dummy  XM_output_mirr_combined_with_dummy_0
timestamp 1662903677
transform 1 0 16600 0 1 14200
box -17600 -7400 35500 15000
use opamp_realcomp3_usefinger  opamp_realcomp3_usefinger_0
timestamp 1662836520
transform 1 0 4380 0 1 -594
box -5380 594 6776 6403
use sky130_fd_pr__nfet_01v8_lvt_E2U6GT  sky130_fd_pr__nfet_01v8_lvt_E2U6GT_0
timestamp 1672431769
transform 1 0 12196 0 1 1359
box -596 -679 596 679
use sky130_fd_pr__nfet_01v8_lvt_H8V8HY  sky130_fd_pr__nfet_01v8_lvt_H8V8HY_0
timestamp 1672431769
transform 1 0 13096 0 1 859
box -396 -1179 396 1179
use sky130_fd_pr__pfet_01v8_lvt_MUVN4U  sky130_fd_pr__pfet_01v8_lvt_MUVN4U_0
timestamp 1672432293
transform 1 0 12412 0 1 2626
box -812 -466 812 466
use sky130_fd_pr__res_high_po_1p41_EL7NMZ  sky130_fd_pr__res_high_po_1p41_EL7NMZ_0
timestamp 1672432498
transform 0 -1 22598 1 0 -733
box -307 -5598 307 5598
use sky130_fd_pr__res_high_po_1p41_G3LFBQ  sky130_fd_pr__res_high_po_1p41_G3LFBQ_0
timestamp 1672432498
transform 0 1 27998 -1 0 -213
box -307 -10998 307 10998
<< labels >>
flabel metal3 13210 4940 13250 5000 0 FreeSans 960 0 0 0 C
flabel space 14620 4940 14660 5000 0 FreeSans 960 0 0 0 C
flabel space 13200 3850 13240 3910 0 FreeSans 960 0 0 0 C
flabel space 14620 3870 14660 3930 0 FreeSans 960 0 0 0 C
flabel metal3 16700 2600 16900 3000 0 FreeSans 1600 0 0 0 vd4
flabel space 16600 21600 16900 21800 0 FreeSans 1600 0 0 0 C
flabel space 16600 14200 16900 14400 0 FreeSans 1600 0 0 0 C
flabel space 34200 14200 34500 14400 0 FreeSans 1600 0 0 0 C
flabel space 34200 21600 34500 21800 0 FreeSans 1600 0 0 0 C
<< end >>
