magic
tech sky130A
timestamp 1671764736
<< pwell >>
rect -1044 -155 1043 155
<< nmoslvt >>
rect -944 -50 -929 50
rect -896 -50 -881 50
rect -848 -50 -833 50
rect -800 -50 -785 50
rect -752 -50 -737 50
rect -704 -50 -689 50
rect -656 -50 -641 50
rect -608 -50 -593 50
rect -560 -50 -545 50
rect -512 -50 -497 50
rect -464 -50 -449 50
rect -416 -50 -401 50
rect -368 -50 -353 50
rect -320 -50 -305 50
rect -272 -50 -257 50
rect -224 -50 -209 50
rect -176 -50 -161 50
rect -128 -50 -113 50
rect -80 -50 -65 50
rect -32 -50 -17 50
rect 16 -50 31 50
rect 64 -50 79 50
rect 112 -50 127 50
rect 160 -50 175 50
rect 208 -50 223 50
rect 256 -50 271 50
rect 304 -50 319 50
rect 352 -50 367 50
rect 400 -50 415 50
rect 448 -50 463 50
rect 496 -50 511 50
rect 544 -50 559 50
rect 592 -50 607 50
rect 640 -50 655 50
rect 688 -50 703 50
rect 736 -50 751 50
rect 784 -50 799 50
rect 832 -50 847 50
rect 880 -50 895 50
rect 928 -50 943 50
<< ndiff >>
rect -975 44 -944 50
rect -975 -44 -969 44
rect -952 -44 -944 44
rect -975 -50 -944 -44
rect -929 44 -896 50
rect -929 -44 -921 44
rect -904 -44 -896 44
rect -929 -50 -896 -44
rect -881 44 -848 50
rect -881 -44 -873 44
rect -856 -44 -848 44
rect -881 -50 -848 -44
rect -833 44 -800 50
rect -833 -44 -825 44
rect -808 -44 -800 44
rect -833 -50 -800 -44
rect -785 44 -752 50
rect -785 -44 -777 44
rect -760 -44 -752 44
rect -785 -50 -752 -44
rect -737 44 -704 50
rect -737 -44 -729 44
rect -712 -44 -704 44
rect -737 -50 -704 -44
rect -689 44 -656 50
rect -689 -44 -681 44
rect -664 -44 -656 44
rect -689 -50 -656 -44
rect -641 44 -608 50
rect -641 -44 -633 44
rect -616 -44 -608 44
rect -641 -50 -608 -44
rect -593 44 -560 50
rect -593 -44 -585 44
rect -568 -44 -560 44
rect -593 -50 -560 -44
rect -545 44 -512 50
rect -545 -44 -537 44
rect -520 -44 -512 44
rect -545 -50 -512 -44
rect -497 44 -464 50
rect -497 -44 -489 44
rect -472 -44 -464 44
rect -497 -50 -464 -44
rect -449 44 -416 50
rect -449 -44 -441 44
rect -424 -44 -416 44
rect -449 -50 -416 -44
rect -401 44 -368 50
rect -401 -44 -393 44
rect -376 -44 -368 44
rect -401 -50 -368 -44
rect -353 44 -320 50
rect -353 -44 -345 44
rect -328 -44 -320 44
rect -353 -50 -320 -44
rect -305 44 -272 50
rect -305 -44 -297 44
rect -280 -44 -272 44
rect -305 -50 -272 -44
rect -257 44 -224 50
rect -257 -44 -249 44
rect -232 -44 -224 44
rect -257 -50 -224 -44
rect -209 44 -176 50
rect -209 -44 -201 44
rect -184 -44 -176 44
rect -209 -50 -176 -44
rect -161 44 -128 50
rect -161 -44 -153 44
rect -136 -44 -128 44
rect -161 -50 -128 -44
rect -113 44 -80 50
rect -113 -44 -105 44
rect -88 -44 -80 44
rect -113 -50 -80 -44
rect -65 44 -32 50
rect -65 -44 -57 44
rect -40 -44 -32 44
rect -65 -50 -32 -44
rect -17 44 16 50
rect -17 -44 -9 44
rect 8 -44 16 44
rect -17 -50 16 -44
rect 31 44 64 50
rect 31 -44 39 44
rect 56 -44 64 44
rect 31 -50 64 -44
rect 79 44 112 50
rect 79 -44 87 44
rect 104 -44 112 44
rect 79 -50 112 -44
rect 127 44 160 50
rect 127 -44 135 44
rect 152 -44 160 44
rect 127 -50 160 -44
rect 175 44 208 50
rect 175 -44 183 44
rect 200 -44 208 44
rect 175 -50 208 -44
rect 223 44 256 50
rect 223 -44 231 44
rect 248 -44 256 44
rect 223 -50 256 -44
rect 271 44 304 50
rect 271 -44 279 44
rect 296 -44 304 44
rect 271 -50 304 -44
rect 319 44 352 50
rect 319 -44 327 44
rect 344 -44 352 44
rect 319 -50 352 -44
rect 367 44 400 50
rect 367 -44 375 44
rect 392 -44 400 44
rect 367 -50 400 -44
rect 415 44 448 50
rect 415 -44 423 44
rect 440 -44 448 44
rect 415 -50 448 -44
rect 463 44 496 50
rect 463 -44 471 44
rect 488 -44 496 44
rect 463 -50 496 -44
rect 511 44 544 50
rect 511 -44 519 44
rect 536 -44 544 44
rect 511 -50 544 -44
rect 559 44 592 50
rect 559 -44 567 44
rect 584 -44 592 44
rect 559 -50 592 -44
rect 607 44 640 50
rect 607 -44 615 44
rect 632 -44 640 44
rect 607 -50 640 -44
rect 655 44 688 50
rect 655 -44 663 44
rect 680 -44 688 44
rect 655 -50 688 -44
rect 703 44 736 50
rect 703 -44 711 44
rect 728 -44 736 44
rect 703 -50 736 -44
rect 751 44 784 50
rect 751 -44 759 44
rect 776 -44 784 44
rect 751 -50 784 -44
rect 799 44 832 50
rect 799 -44 807 44
rect 824 -44 832 44
rect 799 -50 832 -44
rect 847 44 880 50
rect 847 -44 855 44
rect 872 -44 880 44
rect 847 -50 880 -44
rect 895 44 928 50
rect 895 -44 903 44
rect 920 -44 928 44
rect 895 -50 928 -44
rect 943 44 974 50
rect 943 -44 951 44
rect 968 -44 974 44
rect 943 -50 974 -44
<< ndiffc >>
rect -969 -44 -952 44
rect -921 -44 -904 44
rect -873 -44 -856 44
rect -825 -44 -808 44
rect -777 -44 -760 44
rect -729 -44 -712 44
rect -681 -44 -664 44
rect -633 -44 -616 44
rect -585 -44 -568 44
rect -537 -44 -520 44
rect -489 -44 -472 44
rect -441 -44 -424 44
rect -393 -44 -376 44
rect -345 -44 -328 44
rect -297 -44 -280 44
rect -249 -44 -232 44
rect -201 -44 -184 44
rect -153 -44 -136 44
rect -105 -44 -88 44
rect -57 -44 -40 44
rect -9 -44 8 44
rect 39 -44 56 44
rect 87 -44 104 44
rect 135 -44 152 44
rect 183 -44 200 44
rect 231 -44 248 44
rect 279 -44 296 44
rect 327 -44 344 44
rect 375 -44 392 44
rect 423 -44 440 44
rect 471 -44 488 44
rect 519 -44 536 44
rect 567 -44 584 44
rect 615 -44 632 44
rect 663 -44 680 44
rect 711 -44 728 44
rect 759 -44 776 44
rect 807 -44 824 44
rect 855 -44 872 44
rect 903 -44 920 44
rect 951 -44 968 44
<< psubdiff >>
rect -1026 120 -978 137
rect 977 120 1025 137
rect -1026 89 -1009 120
rect 1008 89 1025 120
rect -1026 -120 -1009 -89
rect 1008 -120 1025 -89
rect -1026 -137 -978 -120
rect 977 -137 1025 -120
<< psubdiffcont >>
rect -978 120 977 137
rect -1026 -89 -1009 89
rect 1008 -89 1025 89
rect -978 -137 977 -120
<< poly >>
rect -944 50 -929 63
rect -896 50 -881 63
rect -848 50 -833 63
rect -800 50 -785 63
rect -752 50 -737 63
rect -704 50 -689 63
rect -656 50 -641 63
rect -608 50 -593 63
rect -560 50 -545 63
rect -512 50 -497 63
rect -464 50 -449 63
rect -416 50 -401 63
rect -368 50 -353 63
rect -320 50 -305 63
rect -272 50 -257 63
rect -224 50 -209 63
rect -176 50 -161 63
rect -128 50 -113 63
rect -80 50 -65 63
rect -32 50 -17 63
rect 16 50 31 63
rect 64 50 79 63
rect 112 50 127 63
rect 160 50 175 63
rect 208 50 223 63
rect 256 50 271 63
rect 304 50 319 63
rect 352 50 367 63
rect 400 50 415 63
rect 448 50 463 63
rect 496 50 511 63
rect 544 50 559 63
rect 592 50 607 63
rect 640 50 655 63
rect 688 50 703 63
rect 736 50 751 63
rect 784 50 799 63
rect 832 50 847 63
rect 880 50 895 63
rect 928 50 943 63
rect -944 -61 -929 -50
rect -953 -63 -920 -61
rect -896 -63 -881 -50
rect -848 -61 -833 -50
rect -857 -63 -824 -61
rect -800 -63 -785 -50
rect -752 -61 -737 -50
rect -761 -63 -728 -61
rect -704 -63 -689 -50
rect -656 -61 -641 -50
rect -665 -63 -632 -61
rect -608 -63 -593 -50
rect -560 -61 -545 -50
rect -569 -63 -536 -61
rect -512 -63 -497 -50
rect -464 -61 -449 -50
rect -473 -63 -440 -61
rect -416 -63 -401 -50
rect -368 -61 -353 -50
rect -377 -63 -344 -61
rect -320 -63 -305 -50
rect -272 -61 -257 -50
rect -281 -63 -248 -61
rect -224 -63 -209 -50
rect -176 -61 -161 -50
rect -185 -63 -152 -61
rect -128 -63 -113 -50
rect -80 -61 -65 -50
rect -89 -63 -56 -61
rect -32 -63 -17 -50
rect 16 -61 31 -50
rect 7 -63 40 -61
rect 64 -63 79 -50
rect 112 -61 127 -50
rect 103 -63 136 -61
rect 160 -63 175 -50
rect 208 -61 223 -50
rect 199 -63 232 -61
rect 256 -63 271 -50
rect 304 -61 319 -50
rect 295 -63 328 -61
rect 352 -63 367 -50
rect 400 -61 415 -50
rect 391 -63 424 -61
rect 448 -63 463 -50
rect 496 -61 511 -50
rect 487 -63 520 -61
rect 544 -63 559 -50
rect 592 -61 607 -50
rect 583 -63 616 -61
rect 640 -63 655 -50
rect 688 -61 703 -50
rect 679 -63 712 -61
rect 736 -63 751 -50
rect 784 -61 799 -50
rect 775 -63 808 -61
rect 832 -63 847 -50
rect 880 -61 895 -50
rect 871 -63 904 -61
rect 928 -63 943 -50
rect -953 -69 943 -63
rect -953 -81 15 -69
rect -953 -94 -920 -81
rect -857 -94 -824 -81
rect -761 -94 -728 -81
rect -665 -94 -632 -81
rect -569 -94 -536 -81
rect -473 -94 -440 -81
rect -377 -94 -344 -81
rect -281 -94 -248 -81
rect -185 -94 -152 -81
rect -89 -94 -56 -81
rect 7 -86 15 -81
rect 32 -81 943 -69
rect 32 -86 40 -81
rect 7 -94 40 -86
rect 103 -94 136 -81
rect 199 -94 232 -81
rect 295 -94 328 -81
rect 391 -94 424 -81
rect 487 -94 520 -81
rect 583 -94 616 -81
rect 679 -94 712 -81
rect 775 -94 808 -81
rect 871 -94 904 -81
<< polycont >>
rect 15 -86 32 -69
<< locali >>
rect -1026 120 -978 137
rect 977 120 1025 137
rect -1026 89 -1009 120
rect 1008 89 1025 120
rect -969 44 -952 52
rect -969 -52 -952 -44
rect -921 44 -904 52
rect -921 -52 -904 -44
rect -873 44 -856 52
rect -873 -52 -856 -44
rect -825 44 -808 52
rect -825 -52 -808 -44
rect -777 44 -760 52
rect -777 -52 -760 -44
rect -729 44 -712 52
rect -729 -52 -712 -44
rect -681 44 -664 52
rect -681 -52 -664 -44
rect -633 44 -616 52
rect -633 -52 -616 -44
rect -585 44 -568 52
rect -585 -52 -568 -44
rect -537 44 -520 52
rect -537 -52 -520 -44
rect -489 44 -472 52
rect -489 -52 -472 -44
rect -441 44 -424 52
rect -441 -52 -424 -44
rect -393 44 -376 52
rect -393 -52 -376 -44
rect -345 44 -328 52
rect -345 -52 -328 -44
rect -297 44 -280 52
rect -297 -52 -280 -44
rect -249 44 -232 52
rect -249 -52 -232 -44
rect -201 44 -184 52
rect -201 -52 -184 -44
rect -153 44 -136 52
rect -153 -52 -136 -44
rect -105 44 -88 52
rect -105 -52 -88 -44
rect -57 44 -40 52
rect -57 -52 -40 -44
rect -9 44 8 52
rect -9 -52 8 -44
rect 39 44 56 52
rect 39 -52 56 -44
rect 87 44 104 52
rect 87 -52 104 -44
rect 135 44 152 52
rect 135 -52 152 -44
rect 183 44 200 52
rect 183 -52 200 -44
rect 231 44 248 52
rect 231 -52 248 -44
rect 279 44 296 52
rect 279 -52 296 -44
rect 327 44 344 52
rect 327 -52 344 -44
rect 375 44 392 52
rect 375 -52 392 -44
rect 423 44 440 52
rect 423 -52 440 -44
rect 471 44 488 52
rect 471 -52 488 -44
rect 519 44 536 52
rect 519 -52 536 -44
rect 567 44 584 52
rect 567 -52 584 -44
rect 615 44 632 52
rect 615 -52 632 -44
rect 663 44 680 52
rect 663 -52 680 -44
rect 711 44 728 52
rect 711 -52 728 -44
rect 759 44 776 52
rect 759 -52 776 -44
rect 807 44 824 52
rect 807 -52 824 -44
rect 855 44 872 52
rect 855 -52 872 -44
rect 903 44 920 52
rect 903 -52 920 -44
rect 951 44 968 52
rect 951 -52 968 -44
rect 7 -86 15 -69
rect 32 -86 40 -69
rect -1026 -120 -1009 -89
rect 1008 -120 1025 -89
rect -1026 -137 -978 -120
rect 977 -137 1025 -120
<< viali >>
rect -969 -44 -952 44
rect -921 -44 -904 44
rect -873 -44 -856 44
rect -825 -44 -808 44
rect -777 -44 -760 44
rect -729 -44 -712 44
rect -681 -44 -664 44
rect -633 -44 -616 44
rect -585 -44 -568 44
rect -537 -44 -520 44
rect -489 -44 -472 44
rect -441 -44 -424 44
rect -393 -44 -376 44
rect -345 -44 -328 44
rect -297 -44 -280 44
rect -249 -44 -232 44
rect -201 -44 -184 44
rect -153 -44 -136 44
rect -105 -44 -88 44
rect -57 -44 -40 44
rect -9 -44 8 44
rect 39 -44 56 44
rect 87 -44 104 44
rect 135 -44 152 44
rect 183 -44 200 44
rect 231 -44 248 44
rect 279 -44 296 44
rect 327 -44 344 44
rect 375 -44 392 44
rect 423 -44 440 44
rect 471 -44 488 44
rect 519 -44 536 44
rect 567 -44 584 44
rect 615 -44 632 44
rect 663 -44 680 44
rect 711 -44 728 44
rect 759 -44 776 44
rect 807 -44 824 44
rect 855 -44 872 44
rect 903 -44 920 44
rect 951 -44 968 44
rect 15 -86 32 -69
<< metal1 >>
rect -972 44 -949 50
rect -972 -18 -969 44
rect -977 -21 -969 -18
rect -952 -18 -949 44
rect -929 47 -896 50
rect -929 21 -926 47
rect -899 21 -896 47
rect -929 18 -921 21
rect -952 -21 -944 -18
rect -977 -47 -974 -21
rect -947 -47 -944 -21
rect -977 -50 -944 -47
rect -924 -44 -921 18
rect -904 18 -896 21
rect -876 44 -853 50
rect -904 -44 -901 18
rect -876 -18 -873 44
rect -924 -50 -901 -44
rect -881 -21 -873 -18
rect -856 -18 -853 44
rect -833 47 -800 50
rect -833 21 -830 47
rect -803 21 -800 47
rect -833 18 -825 21
rect -856 -21 -848 -18
rect -881 -47 -878 -21
rect -851 -47 -848 -21
rect -881 -50 -848 -47
rect -828 -44 -825 18
rect -808 18 -800 21
rect -780 44 -757 50
rect -808 -44 -805 18
rect -780 -18 -777 44
rect -828 -50 -805 -44
rect -785 -21 -777 -18
rect -760 -18 -757 44
rect -737 47 -704 50
rect -737 21 -734 47
rect -707 21 -704 47
rect -737 18 -729 21
rect -760 -21 -752 -18
rect -785 -47 -782 -21
rect -755 -47 -752 -21
rect -785 -50 -752 -47
rect -732 -44 -729 18
rect -712 18 -704 21
rect -684 44 -661 50
rect -712 -44 -709 18
rect -684 -18 -681 44
rect -732 -50 -709 -44
rect -689 -21 -681 -18
rect -664 -18 -661 44
rect -641 47 -608 50
rect -641 21 -638 47
rect -611 21 -608 47
rect -641 18 -633 21
rect -664 -21 -656 -18
rect -689 -47 -686 -21
rect -659 -47 -656 -21
rect -689 -50 -656 -47
rect -636 -44 -633 18
rect -616 18 -608 21
rect -588 44 -565 50
rect -616 -44 -613 18
rect -588 -18 -585 44
rect -636 -50 -613 -44
rect -593 -21 -585 -18
rect -568 -18 -565 44
rect -545 47 -512 50
rect -545 21 -542 47
rect -515 21 -512 47
rect -545 18 -537 21
rect -568 -21 -560 -18
rect -593 -47 -590 -21
rect -563 -47 -560 -21
rect -593 -50 -560 -47
rect -540 -44 -537 18
rect -520 18 -512 21
rect -492 44 -469 50
rect -520 -44 -517 18
rect -492 -18 -489 44
rect -540 -50 -517 -44
rect -497 -21 -489 -18
rect -472 -18 -469 44
rect -449 47 -416 50
rect -449 21 -446 47
rect -419 21 -416 47
rect -449 18 -441 21
rect -472 -21 -464 -18
rect -497 -47 -494 -21
rect -467 -47 -464 -21
rect -497 -50 -464 -47
rect -444 -44 -441 18
rect -424 18 -416 21
rect -396 44 -373 50
rect -424 -44 -421 18
rect -396 -18 -393 44
rect -444 -50 -421 -44
rect -401 -21 -393 -18
rect -376 -18 -373 44
rect -353 47 -320 50
rect -353 21 -350 47
rect -323 21 -320 47
rect -353 18 -345 21
rect -376 -21 -368 -18
rect -401 -47 -398 -21
rect -371 -47 -368 -21
rect -401 -50 -368 -47
rect -348 -44 -345 18
rect -328 18 -320 21
rect -300 44 -277 50
rect -328 -44 -325 18
rect -300 -18 -297 44
rect -348 -50 -325 -44
rect -305 -21 -297 -18
rect -280 -18 -277 44
rect -257 47 -224 50
rect -257 21 -254 47
rect -227 21 -224 47
rect -257 18 -249 21
rect -280 -21 -272 -18
rect -305 -47 -302 -21
rect -275 -47 -272 -21
rect -305 -50 -272 -47
rect -252 -44 -249 18
rect -232 18 -224 21
rect -204 44 -181 50
rect -232 -44 -229 18
rect -204 -18 -201 44
rect -252 -50 -229 -44
rect -209 -21 -201 -18
rect -184 -18 -181 44
rect -161 47 -128 50
rect -161 21 -158 47
rect -131 21 -128 47
rect -161 18 -153 21
rect -184 -21 -176 -18
rect -209 -47 -206 -21
rect -179 -47 -176 -21
rect -209 -50 -176 -47
rect -156 -44 -153 18
rect -136 18 -128 21
rect -108 44 -85 50
rect -136 -44 -133 18
rect -108 -18 -105 44
rect -156 -50 -133 -44
rect -113 -21 -105 -18
rect -88 -18 -85 44
rect -65 47 -32 50
rect -65 21 -62 47
rect -35 21 -32 47
rect -65 18 -57 21
rect -88 -21 -80 -18
rect -113 -47 -110 -21
rect -83 -47 -80 -21
rect -113 -50 -80 -47
rect -60 -44 -57 18
rect -40 18 -32 21
rect -12 44 11 50
rect -40 -44 -37 18
rect -12 -18 -9 44
rect -60 -50 -37 -44
rect -17 -21 -9 -18
rect 8 -18 11 44
rect 31 47 64 50
rect 31 21 34 47
rect 61 21 64 47
rect 31 18 39 21
rect 8 -21 16 -18
rect -17 -47 -14 -21
rect 13 -47 16 -21
rect -17 -50 16 -47
rect 36 -44 39 18
rect 56 18 64 21
rect 84 44 107 50
rect 56 -44 59 18
rect 84 -18 87 44
rect 36 -50 59 -44
rect 79 -21 87 -18
rect 104 -18 107 44
rect 127 47 160 50
rect 127 21 130 47
rect 157 21 160 47
rect 127 18 135 21
rect 104 -21 112 -18
rect 79 -47 82 -21
rect 109 -47 112 -21
rect 79 -50 112 -47
rect 132 -44 135 18
rect 152 18 160 21
rect 180 44 203 50
rect 152 -44 155 18
rect 180 -18 183 44
rect 132 -50 155 -44
rect 175 -21 183 -18
rect 200 -18 203 44
rect 223 47 256 50
rect 223 21 226 47
rect 253 21 256 47
rect 223 18 231 21
rect 200 -21 208 -18
rect 175 -47 178 -21
rect 205 -47 208 -21
rect 175 -50 208 -47
rect 228 -44 231 18
rect 248 18 256 21
rect 276 44 299 50
rect 248 -44 251 18
rect 276 -18 279 44
rect 228 -50 251 -44
rect 271 -21 279 -18
rect 296 -18 299 44
rect 319 47 352 50
rect 319 21 322 47
rect 349 21 352 47
rect 319 18 327 21
rect 296 -21 304 -18
rect 271 -47 274 -21
rect 301 -47 304 -21
rect 271 -50 304 -47
rect 324 -44 327 18
rect 344 18 352 21
rect 372 44 395 50
rect 344 -44 347 18
rect 372 -18 375 44
rect 324 -50 347 -44
rect 367 -21 375 -18
rect 392 -18 395 44
rect 415 47 448 50
rect 415 21 418 47
rect 445 21 448 47
rect 415 18 423 21
rect 392 -21 400 -18
rect 367 -47 370 -21
rect 397 -47 400 -21
rect 367 -50 400 -47
rect 420 -44 423 18
rect 440 18 448 21
rect 468 44 491 50
rect 440 -44 443 18
rect 468 -18 471 44
rect 420 -50 443 -44
rect 463 -21 471 -18
rect 488 -18 491 44
rect 511 47 544 50
rect 511 21 514 47
rect 541 21 544 47
rect 511 18 519 21
rect 488 -21 496 -18
rect 463 -47 466 -21
rect 493 -47 496 -21
rect 463 -50 496 -47
rect 516 -44 519 18
rect 536 18 544 21
rect 564 44 587 50
rect 536 -44 539 18
rect 564 -18 567 44
rect 516 -50 539 -44
rect 559 -21 567 -18
rect 584 -18 587 44
rect 607 47 640 50
rect 607 21 610 47
rect 637 21 640 47
rect 607 18 615 21
rect 584 -21 592 -18
rect 559 -47 562 -21
rect 589 -47 592 -21
rect 559 -50 592 -47
rect 612 -44 615 18
rect 632 18 640 21
rect 660 44 683 50
rect 632 -44 635 18
rect 660 -18 663 44
rect 612 -50 635 -44
rect 655 -21 663 -18
rect 680 -18 683 44
rect 703 47 736 50
rect 703 21 706 47
rect 733 21 736 47
rect 703 18 711 21
rect 680 -21 688 -18
rect 655 -47 658 -21
rect 685 -47 688 -21
rect 655 -50 688 -47
rect 708 -44 711 18
rect 728 18 736 21
rect 756 44 779 50
rect 728 -44 731 18
rect 756 -18 759 44
rect 708 -50 731 -44
rect 751 -21 759 -18
rect 776 -18 779 44
rect 799 47 832 50
rect 799 21 802 47
rect 829 21 832 47
rect 799 18 807 21
rect 776 -21 784 -18
rect 751 -47 754 -21
rect 781 -47 784 -21
rect 751 -50 784 -47
rect 804 -44 807 18
rect 824 18 832 21
rect 852 44 875 50
rect 824 -44 827 18
rect 852 -18 855 44
rect 804 -50 827 -44
rect 847 -21 855 -18
rect 872 -18 875 44
rect 895 47 928 50
rect 895 21 898 47
rect 925 21 928 47
rect 895 18 903 21
rect 872 -21 880 -18
rect 847 -47 850 -21
rect 877 -47 880 -21
rect 847 -50 880 -47
rect 900 -44 903 18
rect 920 18 928 21
rect 948 44 971 50
rect 920 -44 923 18
rect 948 -18 951 44
rect 900 -50 923 -44
rect 943 -21 951 -18
rect 968 -18 971 44
rect 968 -21 976 -18
rect 943 -47 946 -21
rect 973 -47 976 -21
rect 943 -50 976 -47
rect -954 -69 943 -66
rect -954 -86 15 -69
rect 32 -86 943 -69
rect -954 -89 943 -86
<< via1 >>
rect -926 44 -899 47
rect -926 21 -921 44
rect -921 21 -904 44
rect -904 21 -899 44
rect -974 -44 -969 -21
rect -969 -44 -952 -21
rect -952 -44 -947 -21
rect -974 -47 -947 -44
rect -830 44 -803 47
rect -830 21 -825 44
rect -825 21 -808 44
rect -808 21 -803 44
rect -878 -44 -873 -21
rect -873 -44 -856 -21
rect -856 -44 -851 -21
rect -878 -47 -851 -44
rect -734 44 -707 47
rect -734 21 -729 44
rect -729 21 -712 44
rect -712 21 -707 44
rect -782 -44 -777 -21
rect -777 -44 -760 -21
rect -760 -44 -755 -21
rect -782 -47 -755 -44
rect -638 44 -611 47
rect -638 21 -633 44
rect -633 21 -616 44
rect -616 21 -611 44
rect -686 -44 -681 -21
rect -681 -44 -664 -21
rect -664 -44 -659 -21
rect -686 -47 -659 -44
rect -542 44 -515 47
rect -542 21 -537 44
rect -537 21 -520 44
rect -520 21 -515 44
rect -590 -44 -585 -21
rect -585 -44 -568 -21
rect -568 -44 -563 -21
rect -590 -47 -563 -44
rect -446 44 -419 47
rect -446 21 -441 44
rect -441 21 -424 44
rect -424 21 -419 44
rect -494 -44 -489 -21
rect -489 -44 -472 -21
rect -472 -44 -467 -21
rect -494 -47 -467 -44
rect -350 44 -323 47
rect -350 21 -345 44
rect -345 21 -328 44
rect -328 21 -323 44
rect -398 -44 -393 -21
rect -393 -44 -376 -21
rect -376 -44 -371 -21
rect -398 -47 -371 -44
rect -254 44 -227 47
rect -254 21 -249 44
rect -249 21 -232 44
rect -232 21 -227 44
rect -302 -44 -297 -21
rect -297 -44 -280 -21
rect -280 -44 -275 -21
rect -302 -47 -275 -44
rect -158 44 -131 47
rect -158 21 -153 44
rect -153 21 -136 44
rect -136 21 -131 44
rect -206 -44 -201 -21
rect -201 -44 -184 -21
rect -184 -44 -179 -21
rect -206 -47 -179 -44
rect -62 44 -35 47
rect -62 21 -57 44
rect -57 21 -40 44
rect -40 21 -35 44
rect -110 -44 -105 -21
rect -105 -44 -88 -21
rect -88 -44 -83 -21
rect -110 -47 -83 -44
rect 34 44 61 47
rect 34 21 39 44
rect 39 21 56 44
rect 56 21 61 44
rect -14 -44 -9 -21
rect -9 -44 8 -21
rect 8 -44 13 -21
rect -14 -47 13 -44
rect 130 44 157 47
rect 130 21 135 44
rect 135 21 152 44
rect 152 21 157 44
rect 82 -44 87 -21
rect 87 -44 104 -21
rect 104 -44 109 -21
rect 82 -47 109 -44
rect 226 44 253 47
rect 226 21 231 44
rect 231 21 248 44
rect 248 21 253 44
rect 178 -44 183 -21
rect 183 -44 200 -21
rect 200 -44 205 -21
rect 178 -47 205 -44
rect 322 44 349 47
rect 322 21 327 44
rect 327 21 344 44
rect 344 21 349 44
rect 274 -44 279 -21
rect 279 -44 296 -21
rect 296 -44 301 -21
rect 274 -47 301 -44
rect 418 44 445 47
rect 418 21 423 44
rect 423 21 440 44
rect 440 21 445 44
rect 370 -44 375 -21
rect 375 -44 392 -21
rect 392 -44 397 -21
rect 370 -47 397 -44
rect 514 44 541 47
rect 514 21 519 44
rect 519 21 536 44
rect 536 21 541 44
rect 466 -44 471 -21
rect 471 -44 488 -21
rect 488 -44 493 -21
rect 466 -47 493 -44
rect 610 44 637 47
rect 610 21 615 44
rect 615 21 632 44
rect 632 21 637 44
rect 562 -44 567 -21
rect 567 -44 584 -21
rect 584 -44 589 -21
rect 562 -47 589 -44
rect 706 44 733 47
rect 706 21 711 44
rect 711 21 728 44
rect 728 21 733 44
rect 658 -44 663 -21
rect 663 -44 680 -21
rect 680 -44 685 -21
rect 658 -47 685 -44
rect 802 44 829 47
rect 802 21 807 44
rect 807 21 824 44
rect 824 21 829 44
rect 754 -44 759 -21
rect 759 -44 776 -21
rect 776 -44 781 -21
rect 754 -47 781 -44
rect 898 44 925 47
rect 898 21 903 44
rect 903 21 920 44
rect 920 21 925 44
rect 850 -44 855 -21
rect 855 -44 872 -21
rect 872 -44 877 -21
rect 850 -47 877 -44
rect 946 -44 951 -21
rect 951 -44 968 -21
rect 968 -44 973 -21
rect 946 -47 973 -44
<< metal2 >>
rect -977 84 976 94
rect -977 30 -964 84
rect -862 47 976 84
rect -862 30 -830 47
rect -977 21 -926 30
rect -899 21 -830 30
rect -803 21 -734 47
rect -707 21 -638 47
rect -611 21 -542 47
rect -515 21 -446 47
rect -419 21 -350 47
rect -323 21 -254 47
rect -227 21 -158 47
rect -131 21 -62 47
rect -35 21 34 47
rect 61 21 130 47
rect 157 21 226 47
rect 253 21 322 47
rect 349 21 418 47
rect 445 21 514 47
rect 541 21 610 47
rect 637 21 706 47
rect 733 21 802 47
rect 829 21 898 47
rect 925 21 976 47
rect -977 18 976 21
rect -977 -21 976 -18
rect -977 -47 -974 -21
rect -947 -47 -878 -21
rect -851 -47 -782 -21
rect -755 -47 -686 -21
rect -659 -47 -590 -21
rect -563 -47 -494 -21
rect -467 -47 -398 -21
rect -371 -47 -302 -21
rect -275 -47 -206 -21
rect -179 -47 -110 -21
rect -83 -47 -14 -21
rect 13 -47 82 -21
rect 109 -47 178 -21
rect 205 -47 274 -21
rect 301 -47 370 -21
rect 397 -47 466 -21
rect 493 -47 562 -21
rect 589 -47 658 -21
rect 685 -47 754 -21
rect 781 -47 850 -21
rect 877 -28 946 -21
rect 973 -47 976 -21
rect -977 -85 858 -47
rect 961 -85 976 -47
rect -977 -94 976 -85
<< via2 >>
rect -964 47 -862 84
rect -964 30 -926 47
rect -926 30 -899 47
rect -899 30 -862 47
rect 858 -47 877 -28
rect 877 -47 946 -28
rect 946 -47 961 -28
rect 858 -85 961 -47
<< metal3 >>
rect -977 84 -848 94
rect -977 30 -964 84
rect -862 30 -848 84
rect -977 18 -848 30
rect 847 -28 976 -18
rect 847 -85 858 -28
rect 961 -85 976 -28
rect 847 -94 976 -85
<< properties >>
string FIXED_BBOX -1017 -128 1017 128
string gencell sky130_fd_pr__nfet_01v8_lvt
string library sky130
string parameters w 1.0 l 0.15 m 1 nf 40 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
