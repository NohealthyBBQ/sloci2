magic
tech sky130A
magscale 1 2
timestamp 1672439470
<< locali >>
rect 13564 7094 14704 7128
rect 8418 6908 8862 6946
rect 8792 6570 8876 6584
rect 8792 6480 8810 6570
rect 8862 6480 8876 6570
rect 8792 6462 8876 6480
<< viali >>
rect 8810 6480 8862 6570
<< metal1 >>
rect 8092 7330 8894 7390
rect 8164 7294 8222 7330
rect 13338 7008 13404 7114
rect 13460 7008 14084 7064
rect 8792 6570 8992 6628
rect 8792 6480 8810 6570
rect 8862 6480 8992 6570
rect 8792 6462 8992 6480
<< metal2 >>
rect 12570 7418 13528 7436
rect 7896 7220 8032 7296
rect 12570 7238 13114 7418
rect 13504 7238 13528 7418
rect 12570 7224 13528 7238
rect 8016 6670 8134 7162
rect 12538 7128 13496 7168
rect 12180 7026 13496 7128
rect 12182 6808 13496 7026
rect 8016 6348 8944 6670
rect 10328 5330 10688 6402
rect 10328 4752 10348 5330
rect 10672 4752 10688 5330
rect 10328 4730 10688 4752
<< via2 >>
rect 13114 7238 13504 7418
rect 10348 4752 10672 5330
<< metal3 >>
rect 13092 10162 16584 10562
rect 13102 7418 13528 10162
rect 13102 7238 13114 7418
rect 13504 7238 13528 7418
rect 13102 7224 13528 7238
rect 10328 5330 10690 5348
rect 10328 4752 10348 5330
rect 10672 4752 10690 5330
rect 10328 4730 10690 4752
rect 16084 4118 16894 4590
rect 15256 3866 16200 3932
rect 15256 3658 15372 3866
rect 16130 3658 16200 3866
rect 15256 3528 16200 3658
rect 16442 3878 17386 3952
rect 16442 3670 16488 3878
rect 17246 3670 17386 3878
rect 16442 3548 17386 3670
<< via3 >>
rect 10348 4752 10672 5330
rect 15372 3658 16130 3866
rect 16488 3670 17246 3878
<< metal4 >>
rect 15770 8100 16172 10044
rect 16444 8100 16846 10044
rect 10328 5330 10690 5348
rect 10328 4752 10348 5330
rect 10672 4752 10690 5330
rect 10328 4730 10690 4752
rect 15770 3902 16174 6406
rect 16444 4544 16844 6366
rect 16444 3910 16848 4544
rect 15338 3866 16176 3902
rect 15338 3658 15372 3866
rect 16130 3658 16176 3866
rect 15338 3640 16176 3658
rect 16444 3878 17282 3910
rect 16444 3670 16488 3878
rect 17246 3670 17282 3878
rect 16444 3648 17282 3670
<< via4 >>
rect 10358 4768 10658 5322
<< metal5 >>
rect 10680 4728 10684 5246
use sky130_fd_pr__pfet_01v8_lvt_4Q3NH3  XM1
timestamp 1672093385
transform 1 0 8194 0 1 7192
box -296 -320 294 318
use sky130_fd_pr__pfet_01v8_lvt_SUM7J6  XM2
timestamp 1672092821
transform 1 0 10564 0 -1 6964
box -1768 -538 1766 614
use sky130_fd_pr__nfet_01v8_lvt_J2SMEF  XM3
timestamp 1672090903
transform 1 0 13036 0 1 7196
box -600 -310 598 310
use cap_bank3  cap_bank3_0
timestamp 1672090405
transform -1 0 30718 0 -1 -388
box 4978 -4056 23903 -62
use oscillator_core  oscillator_core_0
timestamp 1672439470
transform 1 0 8824 0 1 6360
box 1504 -1790 14070 3860
<< labels >>
flabel space 16444 7780 16846 10044 1 FreeSans 1600 90 0 0 VCO-OUT2
flabel space 15770 7380 16172 10044 1 FreeSans 1600 90 0 0 VCO-OUT1
flabel space 18104 4728 18456 5540 0 FreeSans 1600 0 0 0 VDD
flabel space 10328 4728 10680 5528 0 FreeSans 1600 0 0 0 VDD
flabel space 7896 7220 8166 7296 0 FreeSans 1600 0 0 0 BIAS
<< end >>
