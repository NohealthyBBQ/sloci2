magic
tech sky130A
magscale 1 2
timestamp 1671746277
<< metal3 >>
rect -750 -500 749 500
<< mimcap >>
rect -650 360 550 400
rect -650 -360 -610 360
rect 510 -360 550 360
rect -650 -400 550 -360
<< mimcapcontact >>
rect -610 -360 510 360
<< metal4 >>
rect -611 360 511 361
rect -611 -360 -610 360
rect 510 -360 511 360
rect -611 -361 511 -360
<< properties >>
string FIXED_BBOX -750 -500 650 500
string gencell sky130_fd_pr__cap_mim_m3_1
string library sky130
string parameters w 6.0 l 4.0 val 51.8 carea 2.00 cperi 0.19 nx 1 ny 1 dummy 0 square 0 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 1 tconnect 1 ccov 100
<< end >>
