* NGSPICE file created from user_analog_project_wrapper.ext - technology: sky130A

.subckt sky130_fd_pr__nfet_01v8_lvt_WKNS5B a_n250_n90# a_n280_n120# a_n342_n90# VSUBS
X0 a_n342_n90# a_n280_n120# a_n250_n90# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=1.3e+12p pd=1.06e+07u as=1.3e+12p ps=1.06e+07u w=1e+06u l=150000u
X1 a_n250_n90# a_n280_n120# a_n342_n90# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 a_n250_n90# a_n280_n120# a_n342_n90# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 a_n342_n90# a_n280_n120# a_n250_n90# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 a_n250_n90# a_n280_n120# a_n342_n90# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 a_n250_n90# a_n280_n120# a_n342_n90# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 a_n342_n90# a_n280_n120# a_n250_n90# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
.ends

.subckt sky130_fd_pr__nfet_01v8_lvt_YTLFGX#0 a_n946_n188# a_n1092_n274# a_n990_n100#
+ a_n898_n100#
X0 a_n898_n100# a_n946_n188# a_n990_n100# a_n1092_n274# sky130_fd_pr__nfet_01v8_lvt ad=3.3e+12p pd=2.66e+07u as=3.59e+12p ps=2.918e+07u w=1e+06u l=150000u
X1 a_n898_n100# a_n946_n188# a_n990_n100# a_n1092_n274# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 a_n990_n100# a_n946_n188# a_n898_n100# a_n1092_n274# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 a_n898_n100# a_n946_n188# a_n990_n100# a_n1092_n274# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 a_n990_n100# a_n946_n188# a_n898_n100# a_n1092_n274# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 a_n898_n100# a_n946_n188# a_n990_n100# a_n1092_n274# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 a_n990_n100# a_n946_n188# a_n898_n100# a_n1092_n274# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 a_n990_n100# a_n946_n188# a_n898_n100# a_n1092_n274# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 a_n898_n100# a_n946_n188# a_n990_n100# a_n1092_n274# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 a_n990_n100# a_n946_n188# a_n898_n100# a_n1092_n274# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10 a_n898_n100# a_n946_n188# a_n990_n100# a_n1092_n274# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11 a_n990_n100# a_n946_n188# a_n898_n100# a_n1092_n274# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12 a_n990_n100# a_n946_n188# a_n898_n100# a_n1092_n274# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13 a_n898_n100# a_n946_n188# a_n990_n100# a_n1092_n274# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X14 a_n990_n100# a_n946_n188# a_n898_n100# a_n1092_n274# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X15 a_n898_n100# a_n946_n188# a_n990_n100# a_n1092_n274# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X16 a_n898_n100# a_n946_n188# a_n990_n100# a_n1092_n274# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X17 a_n990_n100# a_n946_n188# a_n898_n100# a_n1092_n274# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X18 a_n990_n100# a_n946_n188# a_n898_n100# a_n1092_n274# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X19 a_n898_n100# a_n946_n188# a_n990_n100# a_n1092_n274# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
.ends

.subckt oscillator_core m1_7086_2470# VSS cap2 cap1
XXM12 m2_5320_n1360# cap1 cap2 VSS sky130_fd_pr__nfet_01v8_lvt_WKNS5B
XXM23 m1_7086_2470# VSS m2_5320_n1360# VSS sky130_fd_pr__nfet_01v8_lvt_YTLFGX#0
XXM25 m1_7086_2470# VSS m2_5320_n1360# VSS sky130_fd_pr__nfet_01v8_lvt_YTLFGX#0
XXM13 cap2 cap1 m2_5320_n1360# VSS sky130_fd_pr__nfet_01v8_lvt_WKNS5B
XXM14 m2_5320_n1360# cap1 cap2 VSS sky130_fd_pr__nfet_01v8_lvt_WKNS5B
XXM24 m1_7086_2470# VSS m2_5320_n1360# VSS sky130_fd_pr__nfet_01v8_lvt_YTLFGX#0
XXM26 m1_7086_2470# VSS m2_5320_n1360# VSS sky130_fd_pr__nfet_01v8_lvt_YTLFGX#0
XXM15 cap2 cap1 m2_5320_n1360# VSS sky130_fd_pr__nfet_01v8_lvt_WKNS5B
XXM16 cap2 cap1 m2_5320_n1360# VSS sky130_fd_pr__nfet_01v8_lvt_WKNS5B
XXM27 m1_7086_2470# VSS m2_5320_n1360# VSS sky130_fd_pr__nfet_01v8_lvt_YTLFGX#0
XXM17 m2_5320_n1360# cap1 cap2 VSS sky130_fd_pr__nfet_01v8_lvt_WKNS5B
XXM28 m1_7086_2470# VSS m2_5320_n1360# VSS sky130_fd_pr__nfet_01v8_lvt_YTLFGX#0
XXM18 cap2 cap1 m2_5320_n1360# VSS sky130_fd_pr__nfet_01v8_lvt_WKNS5B
XXM19 m2_5320_n1360# cap2 cap1 VSS sky130_fd_pr__nfet_01v8_lvt_WKNS5B
XXM1 cap1 cap2 m2_5320_n1360# VSS sky130_fd_pr__nfet_01v8_lvt_WKNS5B
XXM2 m2_5320_n1360# cap2 cap1 VSS sky130_fd_pr__nfet_01v8_lvt_WKNS5B
XXM3 cap1 cap2 m2_5320_n1360# VSS sky130_fd_pr__nfet_01v8_lvt_WKNS5B
XXM4 m2_5320_n1360# cap2 cap1 VSS sky130_fd_pr__nfet_01v8_lvt_WKNS5B
XXM5 cap1 cap2 m2_5320_n1360# VSS sky130_fd_pr__nfet_01v8_lvt_WKNS5B
XXM6 cap1 cap2 m2_5320_n1360# VSS sky130_fd_pr__nfet_01v8_lvt_WKNS5B
Xsky130_fd_pr__nfet_01v8_lvt_WKNS5B_1 cap1 cap2 m2_5320_n1360# VSS sky130_fd_pr__nfet_01v8_lvt_WKNS5B
XXM7 m2_5320_n1360# cap2 cap1 VSS sky130_fd_pr__nfet_01v8_lvt_WKNS5B
XXM8 cap1 cap2 m2_5320_n1360# VSS sky130_fd_pr__nfet_01v8_lvt_WKNS5B
XXM9 m2_5320_n1360# cap1 cap2 VSS sky130_fd_pr__nfet_01v8_lvt_WKNS5B
XXM21 m1_7086_2470# VSS m2_5320_n1360# VSS sky130_fd_pr__nfet_01v8_lvt_YTLFGX#0
XXM10 cap2 cap1 m2_5320_n1360# VSS sky130_fd_pr__nfet_01v8_lvt_WKNS5B
XXM22 m1_7086_2470# VSS m2_5320_n1360# VSS sky130_fd_pr__nfet_01v8_lvt_YTLFGX#0
XXM11 cap2 cap1 m2_5320_n1360# VSS sky130_fd_pr__nfet_01v8_lvt_WKNS5B
.ends

.subckt sky130_fd_pr__pfet_01v8_lvt_4Q3NH3 a_n100_n198# a_n30_n101# w_n296_n320# a_n158_n101#
X0 a_n30_n101# a_n100_n198# a_n158_n101# w_n296_n320# sky130_fd_pr__pfet_01v8_lvt ad=2.9e+11p pd=2.58e+06u as=5.8e+11p ps=5.16e+06u w=1e+06u l=350000u
X1 a_n158_n101# a_n100_n198# a_n30_n101# w_n296_n320# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=350000u
.ends

.subckt sky130_fd_pr__nfet_01v8_lvt_YTLFGX a_n946_n188# a_n1092_n274# a_n990_n100#
+ a_n898_n100#
X0 a_n898_n100# a_n946_n188# a_n990_n100# a_n1092_n274# sky130_fd_pr__nfet_01v8_lvt ad=3.3e+12p pd=2.66e+07u as=3.59e+12p ps=2.918e+07u w=1e+06u l=150000u
X1 a_n898_n100# a_n946_n188# a_n990_n100# a_n1092_n274# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 a_n990_n100# a_n946_n188# a_n898_n100# a_n1092_n274# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 a_n898_n100# a_n946_n188# a_n990_n100# a_n1092_n274# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 a_n990_n100# a_n946_n188# a_n898_n100# a_n1092_n274# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 a_n898_n100# a_n946_n188# a_n990_n100# a_n1092_n274# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 a_n990_n100# a_n946_n188# a_n898_n100# a_n1092_n274# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 a_n990_n100# a_n946_n188# a_n898_n100# a_n1092_n274# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 a_n898_n100# a_n946_n188# a_n990_n100# a_n1092_n274# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 a_n990_n100# a_n946_n188# a_n898_n100# a_n1092_n274# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10 a_n898_n100# a_n946_n188# a_n990_n100# a_n1092_n274# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11 a_n990_n100# a_n946_n188# a_n898_n100# a_n1092_n274# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12 a_n990_n100# a_n946_n188# a_n898_n100# a_n1092_n274# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13 a_n898_n100# a_n946_n188# a_n990_n100# a_n1092_n274# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X14 a_n990_n100# a_n946_n188# a_n898_n100# a_n1092_n274# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X15 a_n898_n100# a_n946_n188# a_n990_n100# a_n1092_n274# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X16 a_n898_n100# a_n946_n188# a_n990_n100# a_n1092_n274# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X17 a_n990_n100# a_n946_n188# a_n898_n100# a_n1092_n274# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X18 a_n990_n100# a_n946_n188# a_n898_n100# a_n1092_n274# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X19 a_n898_n100# a_n946_n188# a_n990_n100# a_n1092_n274# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
.ends

.subckt sky130_fd_pr__nfet_01v8_lvt_A33GGX a_n2052_n274# a_n1906_n188# a_n1950_n100#
+ a_n1858_n100#
X0 a_n1858_n100# a_n1906_n188# a_n1950_n100# a_n2052_n274# sky130_fd_pr__nfet_01v8_lvt ad=6.6e+12p pd=5.32e+07u as=6.89e+12p ps=5.578e+07u w=1e+06u l=150000u
X1 a_n1858_n100# a_n1906_n188# a_n1950_n100# a_n2052_n274# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 a_n1950_n100# a_n1906_n188# a_n1858_n100# a_n2052_n274# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 a_n1858_n100# a_n1906_n188# a_n1950_n100# a_n2052_n274# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 a_n1950_n100# a_n1906_n188# a_n1858_n100# a_n2052_n274# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 a_n1950_n100# a_n1906_n188# a_n1858_n100# a_n2052_n274# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 a_n1858_n100# a_n1906_n188# a_n1950_n100# a_n2052_n274# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 a_n1858_n100# a_n1906_n188# a_n1950_n100# a_n2052_n274# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 a_n1950_n100# a_n1906_n188# a_n1858_n100# a_n2052_n274# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 a_n1858_n100# a_n1906_n188# a_n1950_n100# a_n2052_n274# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10 a_n1950_n100# a_n1906_n188# a_n1858_n100# a_n2052_n274# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11 a_n1858_n100# a_n1906_n188# a_n1950_n100# a_n2052_n274# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12 a_n1950_n100# a_n1906_n188# a_n1858_n100# a_n2052_n274# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13 a_n1950_n100# a_n1906_n188# a_n1858_n100# a_n2052_n274# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X14 a_n1858_n100# a_n1906_n188# a_n1950_n100# a_n2052_n274# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X15 a_n1858_n100# a_n1906_n188# a_n1950_n100# a_n2052_n274# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X16 a_n1950_n100# a_n1906_n188# a_n1858_n100# a_n2052_n274# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X17 a_n1950_n100# a_n1906_n188# a_n1858_n100# a_n2052_n274# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X18 a_n1950_n100# a_n1906_n188# a_n1858_n100# a_n2052_n274# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X19 a_n1858_n100# a_n1906_n188# a_n1950_n100# a_n2052_n274# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X20 a_n1858_n100# a_n1906_n188# a_n1950_n100# a_n2052_n274# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X21 a_n1950_n100# a_n1906_n188# a_n1858_n100# a_n2052_n274# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X22 a_n1950_n100# a_n1906_n188# a_n1858_n100# a_n2052_n274# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X23 a_n1858_n100# a_n1906_n188# a_n1950_n100# a_n2052_n274# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X24 a_n1858_n100# a_n1906_n188# a_n1950_n100# a_n2052_n274# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X25 a_n1950_n100# a_n1906_n188# a_n1858_n100# a_n2052_n274# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X26 a_n1858_n100# a_n1906_n188# a_n1950_n100# a_n2052_n274# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X27 a_n1950_n100# a_n1906_n188# a_n1858_n100# a_n2052_n274# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X28 a_n1950_n100# a_n1906_n188# a_n1858_n100# a_n2052_n274# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X29 a_n1858_n100# a_n1906_n188# a_n1950_n100# a_n2052_n274# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X30 a_n1950_n100# a_n1906_n188# a_n1858_n100# a_n2052_n274# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X31 a_n1858_n100# a_n1906_n188# a_n1950_n100# a_n2052_n274# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X32 a_n1858_n100# a_n1906_n188# a_n1950_n100# a_n2052_n274# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X33 a_n1950_n100# a_n1906_n188# a_n1858_n100# a_n2052_n274# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X34 a_n1950_n100# a_n1906_n188# a_n1858_n100# a_n2052_n274# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X35 a_n1858_n100# a_n1906_n188# a_n1950_n100# a_n2052_n274# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X36 a_n1858_n100# a_n1906_n188# a_n1950_n100# a_n2052_n274# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X37 a_n1950_n100# a_n1906_n188# a_n1858_n100# a_n2052_n274# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X38 a_n1950_n100# a_n1906_n188# a_n1858_n100# a_n2052_n274# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X39 a_n1858_n100# a_n1906_n188# a_n1950_n100# a_n2052_n274# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
.ends

.subckt sky130_fd_pr__nfet_01v8_lvt_LELFGX a_n2866_n188# a_n3012_n274# a_n2910_n100#
+ a_n2818_n100#
X0 a_n2818_n100# a_n2866_n188# a_n2910_n100# a_n3012_n274# sky130_fd_pr__nfet_01v8_lvt ad=9.9e+12p pd=7.98e+07u as=1.019e+13p ps=8.238e+07u w=1e+06u l=150000u
X1 a_n2818_n100# a_n2866_n188# a_n2910_n100# a_n3012_n274# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 a_n2910_n100# a_n2866_n188# a_n2818_n100# a_n3012_n274# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 a_n2818_n100# a_n2866_n188# a_n2910_n100# a_n3012_n274# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 a_n2910_n100# a_n2866_n188# a_n2818_n100# a_n3012_n274# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 a_n2910_n100# a_n2866_n188# a_n2818_n100# a_n3012_n274# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 a_n2818_n100# a_n2866_n188# a_n2910_n100# a_n3012_n274# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 a_n2818_n100# a_n2866_n188# a_n2910_n100# a_n3012_n274# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 a_n2910_n100# a_n2866_n188# a_n2818_n100# a_n3012_n274# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 a_n2818_n100# a_n2866_n188# a_n2910_n100# a_n3012_n274# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10 a_n2910_n100# a_n2866_n188# a_n2818_n100# a_n3012_n274# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11 a_n2818_n100# a_n2866_n188# a_n2910_n100# a_n3012_n274# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12 a_n2910_n100# a_n2866_n188# a_n2818_n100# a_n3012_n274# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13 a_n2910_n100# a_n2866_n188# a_n2818_n100# a_n3012_n274# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X14 a_n2818_n100# a_n2866_n188# a_n2910_n100# a_n3012_n274# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X15 a_n2910_n100# a_n2866_n188# a_n2818_n100# a_n3012_n274# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X16 a_n2910_n100# a_n2866_n188# a_n2818_n100# a_n3012_n274# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X17 a_n2818_n100# a_n2866_n188# a_n2910_n100# a_n3012_n274# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X18 a_n2818_n100# a_n2866_n188# a_n2910_n100# a_n3012_n274# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X19 a_n2910_n100# a_n2866_n188# a_n2818_n100# a_n3012_n274# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X20 a_n2910_n100# a_n2866_n188# a_n2818_n100# a_n3012_n274# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X21 a_n2818_n100# a_n2866_n188# a_n2910_n100# a_n3012_n274# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X22 a_n2818_n100# a_n2866_n188# a_n2910_n100# a_n3012_n274# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X23 a_n2910_n100# a_n2866_n188# a_n2818_n100# a_n3012_n274# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X24 a_n2818_n100# a_n2866_n188# a_n2910_n100# a_n3012_n274# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X25 a_n2910_n100# a_n2866_n188# a_n2818_n100# a_n3012_n274# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X26 a_n2910_n100# a_n2866_n188# a_n2818_n100# a_n3012_n274# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X27 a_n2910_n100# a_n2866_n188# a_n2818_n100# a_n3012_n274# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X28 a_n2818_n100# a_n2866_n188# a_n2910_n100# a_n3012_n274# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X29 a_n2818_n100# a_n2866_n188# a_n2910_n100# a_n3012_n274# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X30 a_n2910_n100# a_n2866_n188# a_n2818_n100# a_n3012_n274# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X31 a_n2910_n100# a_n2866_n188# a_n2818_n100# a_n3012_n274# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X32 a_n2818_n100# a_n2866_n188# a_n2910_n100# a_n3012_n274# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X33 a_n2818_n100# a_n2866_n188# a_n2910_n100# a_n3012_n274# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X34 a_n2818_n100# a_n2866_n188# a_n2910_n100# a_n3012_n274# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X35 a_n2910_n100# a_n2866_n188# a_n2818_n100# a_n3012_n274# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X36 a_n2818_n100# a_n2866_n188# a_n2910_n100# a_n3012_n274# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X37 a_n2910_n100# a_n2866_n188# a_n2818_n100# a_n3012_n274# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X38 a_n2818_n100# a_n2866_n188# a_n2910_n100# a_n3012_n274# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X39 a_n2818_n100# a_n2866_n188# a_n2910_n100# a_n3012_n274# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X40 a_n2910_n100# a_n2866_n188# a_n2818_n100# a_n3012_n274# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X41 a_n2910_n100# a_n2866_n188# a_n2818_n100# a_n3012_n274# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X42 a_n2818_n100# a_n2866_n188# a_n2910_n100# a_n3012_n274# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X43 a_n2818_n100# a_n2866_n188# a_n2910_n100# a_n3012_n274# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X44 a_n2910_n100# a_n2866_n188# a_n2818_n100# a_n3012_n274# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X45 a_n2818_n100# a_n2866_n188# a_n2910_n100# a_n3012_n274# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X46 a_n2910_n100# a_n2866_n188# a_n2818_n100# a_n3012_n274# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X47 a_n2910_n100# a_n2866_n188# a_n2818_n100# a_n3012_n274# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X48 a_n2818_n100# a_n2866_n188# a_n2910_n100# a_n3012_n274# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X49 a_n2910_n100# a_n2866_n188# a_n2818_n100# a_n3012_n274# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X50 a_n2818_n100# a_n2866_n188# a_n2910_n100# a_n3012_n274# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X51 a_n2818_n100# a_n2866_n188# a_n2910_n100# a_n3012_n274# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X52 a_n2910_n100# a_n2866_n188# a_n2818_n100# a_n3012_n274# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X53 a_n2910_n100# a_n2866_n188# a_n2818_n100# a_n3012_n274# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X54 a_n2910_n100# a_n2866_n188# a_n2818_n100# a_n3012_n274# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X55 a_n2818_n100# a_n2866_n188# a_n2910_n100# a_n3012_n274# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X56 a_n2818_n100# a_n2866_n188# a_n2910_n100# a_n3012_n274# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X57 a_n2910_n100# a_n2866_n188# a_n2818_n100# a_n3012_n274# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X58 a_n2910_n100# a_n2866_n188# a_n2818_n100# a_n3012_n274# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X59 a_n2818_n100# a_n2866_n188# a_n2910_n100# a_n3012_n274# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
.ends

.subckt sky130_fd_pr__nfet_01v8_lvt_648S5X a_n74_n100# a_14_n100# a_n34_n188# a_n176_n274#
X0 a_14_n100# a_n34_n188# a_n74_n100# a_n176_n274# sky130_fd_pr__nfet_01v8_lvt ad=2.9e+11p pd=2.58e+06u as=2.9e+11p ps=2.58e+06u w=1e+06u l=150000u
.ends

.subckt sky130_fd_pr__nfet_01v8_lvt_DJ7QE5 a_n228_n274# a_n126_n100# a_n64_n126# a_n34_n100#
X0 a_n34_n100# a_n64_n126# a_n126_n100# a_n228_n274# sky130_fd_pr__nfet_01v8_lvt ad=3.3e+11p pd=2.66e+06u as=6.2e+11p ps=5.24e+06u w=1e+06u l=150000u
X1 a_n126_n100# a_n64_n126# a_n34_n100# a_n228_n274# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
.ends

.subckt sky130_fd_pr__cap_mim_m3_1_A6B8BZ c1_n1250_n1600# m3_n1350_n1700#
X0 c1_n1250_n1600# m3_n1350_n1700# sky130_fd_pr__cap_mim_m3_1 l=1.6e+07u w=1.2e+07u
.ends

.subckt sky130_fd_pr__nfet_01v8_lvt_HNLS5R a_n324_n274# a_n222_n100# a_n160_n126#
+ a_n130_n100#
X0 a_n130_n100# a_n160_n126# a_n222_n100# a_n324_n274# sky130_fd_pr__nfet_01v8_lvt ad=6.6e+11p pd=5.32e+06u as=9.5e+11p ps=7.9e+06u w=1e+06u l=150000u
X1 a_n222_n100# a_n160_n126# a_n130_n100# a_n324_n274# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 a_n222_n100# a_n160_n126# a_n130_n100# a_n324_n274# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 a_n130_n100# a_n160_n126# a_n222_n100# a_n324_n274# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
.ends

.subckt sky130_fd_pr__nfet_01v8_lvt_B6HS5D a_n318_n100# a_n256_n126# a_n420_n274#
+ a_n226_n100#
X0 a_n226_n100# a_n256_n126# a_n318_n100# a_n420_n274# sky130_fd_pr__nfet_01v8_lvt ad=9.9e+11p pd=7.98e+06u as=1.28e+12p ps=1.056e+07u w=1e+06u l=150000u
X1 a_n318_n100# a_n256_n126# a_n226_n100# a_n420_n274# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 a_n318_n100# a_n256_n126# a_n226_n100# a_n420_n274# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 a_n226_n100# a_n256_n126# a_n318_n100# a_n420_n274# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 a_n226_n100# a_n256_n126# a_n318_n100# a_n420_n274# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 a_n318_n100# a_n256_n126# a_n226_n100# a_n420_n274# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
.ends

.subckt sky130_fd_pr__cap_mim_m3_1_3ZFDVT m3_n450_n500# c1_n350_n400#
X0 c1_n350_n400# m3_n450_n500# sky130_fd_pr__cap_mim_m3_1 l=4e+06u w=3e+06u
.ends

.subckt sky130_fd_pr__cap_mim_m3_1_VCH7EQ c1_n650_n400# m3_n750_n500#
X0 c1_n650_n400# m3_n750_n500# sky130_fd_pr__cap_mim_m3_1 l=4e+06u w=6e+06u
.ends

.subckt sky130_fd_pr__cap_mim_m3_1_MYMY8D c1_n650_n800# m3_n750_n900#
X0 c1_n650_n800# m3_n750_n900# sky130_fd_pr__cap_mim_m3_1 l=8e+06u w=6e+06u
.ends

.subckt sky130_fd_pr__cap_mim_m3_1_CYFFME m3_n1350_n900# c1_n1250_n800#
X0 c1_n1250_n800# m3_n1350_n900# sky130_fd_pr__cap_mim_m3_1 l=8e+06u w=1.2e+07u
.ends

.subckt sky130_fd_pr__nfet_01v8_lvt_9DHFGX a_n612_n274# a_n510_n100# a_n418_n100#
+ a_n466_n188#
X0 a_n510_n100# a_n466_n188# a_n418_n100# a_n612_n274# sky130_fd_pr__nfet_01v8_lvt ad=1.94e+12p pd=1.588e+07u as=1.65e+12p ps=1.33e+07u w=1e+06u l=150000u
X1 a_n418_n100# a_n466_n188# a_n510_n100# a_n612_n274# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 a_n418_n100# a_n466_n188# a_n510_n100# a_n612_n274# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 a_n510_n100# a_n466_n188# a_n418_n100# a_n612_n274# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 a_n510_n100# a_n466_n188# a_n418_n100# a_n612_n274# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 a_n418_n100# a_n466_n188# a_n510_n100# a_n612_n274# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 a_n418_n100# a_n466_n188# a_n510_n100# a_n612_n274# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 a_n510_n100# a_n466_n188# a_n418_n100# a_n612_n274# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 a_n418_n100# a_n466_n188# a_n510_n100# a_n612_n274# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 a_n510_n100# a_n466_n188# a_n418_n100# a_n612_n274# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
.ends

.subckt cap_bank3 m3_14518_n4040# m3_5100_n4040# ctrll5 ctrll4 ctrll2 ctrll3 ctrll1
+ GND
XXM12 ctrll2 GND m2_14442_n2176# m2_12742_n1970# sky130_fd_pr__nfet_01v8_lvt_YTLFGX
XXM13 ctrll3 GND m2_16704_n1564# m2_11726_n1758# sky130_fd_pr__nfet_01v8_lvt_YTLFGX
XXM14 GND ctrll4 m2_18556_n1762# m2_9978_n1770# sky130_fd_pr__nfet_01v8_lvt_A33GGX
XXM15 ctrll5 GND m2_17562_n544# m2_8468_n1256# sky130_fd_pr__nfet_01v8_lvt_LELFGX
XXM1 GND m3_13400_n2830# ctrll1 GND sky130_fd_pr__nfet_01v8_lvt_648S5X
XXM2 GND m2_12742_n1970# ctrll2 GND sky130_fd_pr__nfet_01v8_lvt_DJ7QE5
XXC10 m2_17562_n544# m3_14518_n4040# sky130_fd_pr__cap_mim_m3_1_A6B8BZ
XXM3 GND m2_11726_n1758# ctrll3 GND sky130_fd_pr__nfet_01v8_lvt_HNLS5R
XXM4 GND m2_9978_n1770# ctrll4 GND sky130_fd_pr__nfet_01v8_lvt_HNLS5R
XXM5 GND ctrll5 GND m2_8468_n1256# sky130_fd_pr__nfet_01v8_lvt_B6HS5D
XXM6 GND m3_14648_n2610# ctrll1 GND sky130_fd_pr__nfet_01v8_lvt_648S5X
XXM7 GND m2_14442_n2176# ctrll2 GND sky130_fd_pr__nfet_01v8_lvt_DJ7QE5
XXM9 GND m2_18556_n1762# ctrll4 GND sky130_fd_pr__nfet_01v8_lvt_HNLS5R
XXM8 GND m2_16704_n1564# ctrll3 GND sky130_fd_pr__nfet_01v8_lvt_HNLS5R
XXC1 m3_5100_n4040# m3_13400_n2830# sky130_fd_pr__cap_mim_m3_1_3ZFDVT
XXC2 m2_12742_n1970# m3_5100_n4040# sky130_fd_pr__cap_mim_m3_1_VCH7EQ
XXC3 m2_11726_n1758# m3_5100_n4040# sky130_fd_pr__cap_mim_m3_1_MYMY8D
XXC4 m3_5100_n4040# m2_9978_n1770# sky130_fd_pr__cap_mim_m3_1_CYFFME
XXC5 m2_8468_n1256# m3_5100_n4040# sky130_fd_pr__cap_mim_m3_1_A6B8BZ
XXC7 m2_14442_n2176# m3_14518_n4040# sky130_fd_pr__cap_mim_m3_1_VCH7EQ
XXC6 m3_14518_n4040# m3_14648_n2610# sky130_fd_pr__cap_mim_m3_1_3ZFDVT
XXC8 m2_16704_n1564# m3_14518_n4040# sky130_fd_pr__cap_mim_m3_1_MYMY8D
XXC9 m3_14518_n4040# m2_18556_n1762# sky130_fd_pr__cap_mim_m3_1_CYFFME
XXM10 GND ctrll5 GND m2_17562_n544# sky130_fd_pr__nfet_01v8_lvt_B6HS5D
XXM11 GND m3_13400_n2830# m3_14648_n2610# ctrll1 sky130_fd_pr__nfet_01v8_lvt_9DHFGX
.ends

.subckt sky130_fd_pr__pfet_01v8_lvt_SUM7J6 a_n1502_n319# a_n1680_n432# w_n1768_n538#
+ a_n1630_n319#
X0 a_n1630_n319# a_n1680_n432# a_n1502_n319# w_n1768_n538# sky130_fd_pr__pfet_01v8_lvt ad=7.54e+12p pd=6.708e+07u as=7.54e+12p ps=6.708e+07u w=1e+06u l=350000u
X1 a_n1502_n319# a_n1680_n432# a_n1630_n319# w_n1768_n538# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=350000u
X2 a_n1630_n319# a_n1680_n432# a_n1502_n319# w_n1768_n538# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=350000u
X3 a_n1502_n319# a_n1680_n432# a_n1630_n319# w_n1768_n538# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=350000u
X4 a_n1630_n319# a_n1680_n432# a_n1502_n319# w_n1768_n538# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=350000u
X5 a_n1630_n319# a_n1680_n432# a_n1502_n319# w_n1768_n538# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=350000u
X6 a_n1630_n319# a_n1680_n432# a_n1502_n319# w_n1768_n538# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=350000u
X7 a_n1630_n319# a_n1680_n432# a_n1502_n319# w_n1768_n538# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=350000u
X8 a_n1502_n319# a_n1680_n432# a_n1630_n319# w_n1768_n538# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=350000u
X9 a_n1502_n319# a_n1680_n432# a_n1630_n319# w_n1768_n538# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=350000u
X10 a_n1630_n319# a_n1680_n432# a_n1502_n319# w_n1768_n538# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=350000u
X11 a_n1630_n319# a_n1680_n432# a_n1502_n319# w_n1768_n538# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=350000u
X12 a_n1502_n319# a_n1680_n432# a_n1630_n319# w_n1768_n538# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=350000u
X13 a_n1630_n319# a_n1680_n432# a_n1502_n319# w_n1768_n538# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=350000u
X14 a_n1502_n319# a_n1680_n432# a_n1630_n319# w_n1768_n538# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=350000u
X15 a_n1502_n319# a_n1680_n432# a_n1630_n319# w_n1768_n538# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=350000u
X16 a_n1630_n319# a_n1680_n432# a_n1502_n319# w_n1768_n538# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=350000u
X17 a_n1630_n319# a_n1680_n432# a_n1502_n319# w_n1768_n538# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=350000u
X18 a_n1502_n319# a_n1680_n432# a_n1630_n319# w_n1768_n538# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=350000u
X19 a_n1630_n319# a_n1680_n432# a_n1502_n319# w_n1768_n538# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=350000u
X20 a_n1502_n319# a_n1680_n432# a_n1630_n319# w_n1768_n538# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=350000u
X21 a_n1502_n319# a_n1680_n432# a_n1630_n319# w_n1768_n538# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=350000u
X22 a_n1630_n319# a_n1680_n432# a_n1502_n319# w_n1768_n538# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=350000u
X23 a_n1630_n319# a_n1680_n432# a_n1502_n319# w_n1768_n538# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=350000u
X24 a_n1502_n319# a_n1680_n432# a_n1630_n319# w_n1768_n538# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=350000u
X25 a_n1502_n319# a_n1680_n432# a_n1630_n319# w_n1768_n538# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=350000u
X26 a_n1502_n319# a_n1680_n432# a_n1630_n319# w_n1768_n538# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=350000u
X27 a_n1502_n319# a_n1680_n432# a_n1630_n319# w_n1768_n538# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=350000u
X28 a_n1630_n319# a_n1680_n432# a_n1502_n319# w_n1768_n538# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=350000u
X29 a_n1630_n319# a_n1680_n432# a_n1502_n319# w_n1768_n538# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=350000u
X30 a_n1502_n319# a_n1680_n432# a_n1630_n319# w_n1768_n538# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=350000u
X31 a_n1630_n319# a_n1680_n432# a_n1502_n319# w_n1768_n538# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=350000u
X32 a_n1630_n319# a_n1680_n432# a_n1502_n319# w_n1768_n538# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=350000u
X33 a_n1630_n319# a_n1680_n432# a_n1502_n319# w_n1768_n538# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=350000u
X34 a_n1502_n319# a_n1680_n432# a_n1630_n319# w_n1768_n538# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=350000u
X35 a_n1502_n319# a_n1680_n432# a_n1630_n319# w_n1768_n538# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=350000u
X36 a_n1630_n319# a_n1680_n432# a_n1502_n319# w_n1768_n538# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=350000u
X37 a_n1502_n319# a_n1680_n432# a_n1630_n319# w_n1768_n538# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=350000u
X38 a_n1630_n319# a_n1680_n432# a_n1502_n319# w_n1768_n538# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=350000u
X39 a_n1502_n319# a_n1680_n432# a_n1630_n319# w_n1768_n538# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=350000u
X40 a_n1502_n319# a_n1680_n432# a_n1630_n319# w_n1768_n538# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=350000u
X41 a_n1630_n319# a_n1680_n432# a_n1502_n319# w_n1768_n538# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=350000u
X42 a_n1502_n319# a_n1680_n432# a_n1630_n319# w_n1768_n538# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=350000u
X43 a_n1630_n319# a_n1680_n432# a_n1502_n319# w_n1768_n538# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=350000u
X44 a_n1502_n319# a_n1680_n432# a_n1630_n319# w_n1768_n538# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=350000u
X45 a_n1630_n319# a_n1680_n432# a_n1502_n319# w_n1768_n538# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=350000u
X46 a_n1502_n319# a_n1680_n432# a_n1630_n319# w_n1768_n538# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=350000u
X47 a_n1502_n319# a_n1680_n432# a_n1630_n319# w_n1768_n538# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=350000u
X48 a_n1502_n319# a_n1680_n432# a_n1630_n319# w_n1768_n538# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=350000u
X49 a_n1502_n319# a_n1680_n432# a_n1630_n319# w_n1768_n538# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=350000u
.ends

.subckt sky130_fd_pr__nfet_01v8_lvt_J2SMEF a_n564_n274# a_n418_n172# a_n462_n100#
+ a_n370_n100#
X0 a_n370_n100# a_n418_n172# a_n462_n100# a_n564_n274# sky130_fd_pr__nfet_01v8_lvt ad=1.63e+12p pd=1.326e+07u as=1.63e+12p ps=1.326e+07u w=1e+06u l=150000u
X1 a_n462_n100# a_n418_n172# a_n370_n100# a_n564_n274# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 a_n370_n100# a_n418_n172# a_n462_n100# a_n564_n274# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 a_n462_n100# a_n418_n172# a_n370_n100# a_n564_n274# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 a_n370_n100# a_n418_n172# a_n462_n100# a_n564_n274# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 a_n370_n100# a_n418_n172# a_n462_n100# a_n564_n274# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 a_n462_n100# a_n418_n172# a_n370_n100# a_n564_n274# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 a_n462_n100# a_n418_n172# a_n370_n100# a_n564_n274# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 a_n370_n100# a_n418_n172# a_n462_n100# a_n564_n274# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
.ends

.subckt VCO-assembly cap_bank3_0/ctrll5 cap_bank3_0/ctrll4 cap_bank3_0/ctrll3 cap_bank3_0/ctrll2
+ cap_bank3_0/ctrll1 m2_7896_7220# oscillator_core_0/cap1 oscillator_core_0/cap2 VSUBS
Xoscillator_core_0 m2_12180_7026# VSUBS oscillator_core_0/cap2 oscillator_core_0/cap1
+ oscillator_core
XXM1 m2_7896_7220# m2_7896_7220# oscillator_core_0/cap1 oscillator_core_0/cap1 sky130_fd_pr__pfet_01v8_lvt_4Q3NH3
Xcap_bank3_0 oscillator_core_0/cap1 oscillator_core_0/cap2 cap_bank3_0/ctrll5 cap_bank3_0/ctrll4
+ cap_bank3_0/ctrll2 cap_bank3_0/ctrll3 cap_bank3_0/ctrll1 VSUBS cap_bank3
XXM2 m2_12180_7026# m2_7896_7220# oscillator_core_0/cap1 oscillator_core_0/cap1 sky130_fd_pr__pfet_01v8_lvt_SUM7J6
XXM3 VSUBS m2_12180_7026# m2_12180_7026# VSUBS sky130_fd_pr__nfet_01v8_lvt_J2SMEF
.ends

.subckt sky130_fd_pr__nfet_01v8_lvt_Z6RSN3 a_n1058_n19# a_1000_n19# a_n1160_n193#
+ a_n1000_n107#
X0 a_1000_n19# a_n1000_n107# a_n1058_n19# a_n1160_n193# sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.58e+06u as=1.45e+11p ps=1.58e+06u w=500000u l=1e+07u
.ends

.subckt sky130_fd_pr__res_xhigh_po_5p73_AW8RAB a_n573_5000# a_5637_n5432# a_n8155_n5562#
+ a_5637_5000# a_n5541_5000# a_n1815_n5432# a_n6783_n5432# a_n8025_5000# a_6879_5000#
+ a_n3057_5000# a_n6783_5000# a_3153_n5432# a_n1815_5000# a_n573_n5432# a_n4299_n5432#
+ a_n4299_5000# a_1911_n5432# a_6879_n5432# a_669_n5432# a_n5541_n5432# a_n8025_n5432#
+ a_3153_5000# a_4395_n5432# a_1911_5000# a_669_5000# a_4395_5000# a_n3057_n5432#
X0 a_5637_n5432# a_5637_5000# a_n8155_n5562# sky130_fd_pr__res_xhigh_po_5p73 l=5e+07u
X1 a_n5541_n5432# a_n5541_5000# a_n8155_n5562# sky130_fd_pr__res_xhigh_po_5p73 l=5e+07u
X2 a_1911_n5432# a_1911_5000# a_n8155_n5562# sky130_fd_pr__res_xhigh_po_5p73 l=5e+07u
X3 a_3153_n5432# a_3153_5000# a_n8155_n5562# sky130_fd_pr__res_xhigh_po_5p73 l=5e+07u
X4 a_6879_n5432# a_6879_5000# a_n8155_n5562# sky130_fd_pr__res_xhigh_po_5p73 l=5e+07u
X5 a_n6783_n5432# a_n6783_5000# a_n8155_n5562# sky130_fd_pr__res_xhigh_po_5p73 l=5e+07u
X6 a_n1815_n5432# a_n1815_5000# a_n8155_n5562# sky130_fd_pr__res_xhigh_po_5p73 l=5e+07u
X7 a_4395_n5432# a_4395_5000# a_n8155_n5562# sky130_fd_pr__res_xhigh_po_5p73 l=5e+07u
X8 a_n3057_n5432# a_n3057_5000# a_n8155_n5562# sky130_fd_pr__res_xhigh_po_5p73 l=5e+07u
X9 a_n8025_n5432# a_n8025_5000# a_n8155_n5562# sky130_fd_pr__res_xhigh_po_5p73 l=5e+07u
X10 a_n4299_n5432# a_n4299_5000# a_n8155_n5562# sky130_fd_pr__res_xhigh_po_5p73 l=5e+07u
X11 a_n573_n5432# a_n573_5000# a_n8155_n5562# sky130_fd_pr__res_xhigh_po_5p73 l=5e+07u
X12 a_669_n5432# a_669_5000# a_n8155_n5562# sky130_fd_pr__res_xhigh_po_5p73 l=5e+07u
.ends

.subckt sky130_fd_pr__cap_mim_m3_1_LQXKLG m3_n3150_n12550# c1_n3050_n12450#
X0 c1_n3050_n12450# m3_n3150_n12550# sky130_fd_pr__cap_mim_m3_1 l=3e+07u w=3e+07u
X1 c1_n3050_n12450# m3_n3150_n12550# sky130_fd_pr__cap_mim_m3_1 l=3e+07u w=3e+07u
X2 c1_n3050_n12450# m3_n3150_n12550# sky130_fd_pr__cap_mim_m3_1 l=3e+07u w=3e+07u
X3 c1_n3050_n12450# m3_n3150_n12550# sky130_fd_pr__cap_mim_m3_1 l=3e+07u w=3e+07u
.ends

.subckt rc_model_8cap m1_15830_n15780# VSUBS
Xsky130_fd_pr__nfet_01v8_lvt_Z6RSN3_0 m1_14820_n13900# m1_16920_n14260# VSUBS m1_15830_n15780#
+ sky130_fd_pr__nfet_01v8_lvt_Z6RSN3
Xsky130_fd_pr__nfet_01v8_lvt_Z6RSN3_1 m1_14820_n15340# m1_16920_n14980# VSUBS m1_15830_n15780#
+ sky130_fd_pr__nfet_01v8_lvt_Z6RSN3
Xsky130_fd_pr__nfet_01v8_lvt_Z6RSN3_3 m1_14840_n13120# m1_16920_n13540# VSUBS m1_15830_n15780#
+ sky130_fd_pr__nfet_01v8_lvt_Z6RSN3
Xsky130_fd_pr__nfet_01v8_lvt_Z6RSN3_2 m1_14820_n13900# m1_16920_n13540# VSUBS m1_15830_n15780#
+ sky130_fd_pr__nfet_01v8_lvt_Z6RSN3
Xsky130_fd_pr__nfet_01v8_lvt_Z6RSN3_4 m1_14820_n14620# m1_16920_n14260# VSUBS m1_15830_n15780#
+ sky130_fd_pr__nfet_01v8_lvt_Z6RSN3
Xsky130_fd_pr__nfet_01v8_lvt_Z6RSN3_5 m1_14820_n14620# m1_16920_n14980# VSUBS m1_15830_n15780#
+ sky130_fd_pr__nfet_01v8_lvt_Z6RSN3
Xsky130_fd_pr__nfet_01v8_lvt_Z6RSN3_6 m1_14820_n15340# m1_16920_n15680# VSUBS m1_15830_n15780#
+ sky130_fd_pr__nfet_01v8_lvt_Z6RSN3
Xsky130_fd_pr__nfet_01v8_lvt_Z6RSN3_7 m1_15830_n15780# m1_16920_n15680# VSUBS m1_15830_n15780#
+ sky130_fd_pr__nfet_01v8_lvt_Z6RSN3
Xsky130_fd_pr__res_xhigh_po_5p73_AW8RAB_0 m1_25400_n4800# m1_15000_n11000# VSUBS m1_25400_n12200#
+ m1_25400_400# m1_15000_n3400# m1_15000_1400# VSUBS m1_25400_n12200# m1_25400_n2200#
+ m1_25400_400# m1_15000_n8400# m1_25400_n4800# m1_15000_n6000# m1_15000_n1000# m1_25400_n2200#
+ m1_15000_n8400# m1_14840_n13120# m1_15000_n6000# m1_15000_n1000# m1_15000_1400#
+ m1_25400_n9600# m1_15000_n11000# m1_25400_n7200# m1_25400_n7200# m1_25400_n9600#
+ m1_15000_n3400# sky130_fd_pr__res_xhigh_po_5p73_AW8RAB
Xsky130_fd_pr__cap_mim_m3_1_LQXKLG_0 VSUBS m1_15830_n15780# sky130_fd_pr__cap_mim_m3_1_LQXKLG
Xsky130_fd_pr__cap_mim_m3_1_LQXKLG_1 VSUBS m1_15830_n15780# sky130_fd_pr__cap_mim_m3_1_LQXKLG
.ends

.subckt sky130_fd_pr__nfet_01v8_lvt_WSE2Y6 a_50_n200# a_n108_n200# a_n50_n288# a_n210_n374#
X0 a_50_n200# a_n50_n288# a_n108_n200# a_n210_n374# sky130_fd_pr__nfet_01v8_lvt ad=5.8e+11p pd=4.58e+06u as=5.8e+11p ps=4.58e+06u w=2e+06u l=500000u
.ends

.subckt sky130_fd_pr__pfet_01v8_LDYTSD a_n50_n297# a_50_n200# a_n108_n200# w_n246_n419#
X0 a_50_n200# a_n50_n297# a_n108_n200# w_n246_n419# sky130_fd_pr__pfet_01v8 ad=5.8e+11p pd=4.58e+06u as=5.8e+11p ps=4.58e+06u w=2e+06u l=500000u
.ends

.subckt x3T Vout rst_b pd_in VDD row_sel VSS
Xsky130_fd_pr__nfet_01v8_lvt_WSE2Y6_0 m1_170_n680# Vout row_sel VSS sky130_fd_pr__nfet_01v8_lvt_WSE2Y6
Xsky130_fd_pr__nfet_01v8_lvt_WSE2Y6_1 m1_170_n680# VDD pd_in VSS sky130_fd_pr__nfet_01v8_lvt_WSE2Y6
Xsky130_fd_pr__pfet_01v8_LDYTSD_0 rst_b pd_in VDD VDD sky130_fd_pr__pfet_01v8_LDYTSD
Xsky130_fd_pr__nfet_01v8_lvt_WSE2Y6_2 m1_170_n680# VDD pd_in VSS sky130_fd_pr__nfet_01v8_lvt_WSE2Y6
.ends

.subckt rc_model_4cap m1_15830_n15780# VSUBS
Xsky130_fd_pr__nfet_01v8_lvt_Z6RSN3_0 m1_14820_n13900# m1_16920_n14260# VSUBS m1_15830_n15780#
+ sky130_fd_pr__nfet_01v8_lvt_Z6RSN3
Xsky130_fd_pr__nfet_01v8_lvt_Z6RSN3_1 m1_14820_n15340# m1_16920_n14980# VSUBS m1_15830_n15780#
+ sky130_fd_pr__nfet_01v8_lvt_Z6RSN3
Xsky130_fd_pr__nfet_01v8_lvt_Z6RSN3_3 m1_14840_n13120# m1_16920_n13540# VSUBS m1_15830_n15780#
+ sky130_fd_pr__nfet_01v8_lvt_Z6RSN3
Xsky130_fd_pr__nfet_01v8_lvt_Z6RSN3_2 m1_14820_n13900# m1_16920_n13540# VSUBS m1_15830_n15780#
+ sky130_fd_pr__nfet_01v8_lvt_Z6RSN3
Xsky130_fd_pr__nfet_01v8_lvt_Z6RSN3_4 m1_14820_n14620# m1_16920_n14260# VSUBS m1_15830_n15780#
+ sky130_fd_pr__nfet_01v8_lvt_Z6RSN3
Xsky130_fd_pr__nfet_01v8_lvt_Z6RSN3_5 m1_14820_n14620# m1_16920_n14980# VSUBS m1_15830_n15780#
+ sky130_fd_pr__nfet_01v8_lvt_Z6RSN3
Xsky130_fd_pr__nfet_01v8_lvt_Z6RSN3_6 m1_14820_n15340# m1_16920_n15680# VSUBS m1_15830_n15780#
+ sky130_fd_pr__nfet_01v8_lvt_Z6RSN3
Xsky130_fd_pr__nfet_01v8_lvt_Z6RSN3_7 m1_15830_n15780# m1_16920_n15680# VSUBS m1_15830_n15780#
+ sky130_fd_pr__nfet_01v8_lvt_Z6RSN3
Xsky130_fd_pr__res_xhigh_po_5p73_AW8RAB_0 m1_25400_n4800# m1_15000_n11000# VSUBS m1_25400_n12200#
+ m1_25400_400# m1_15000_n3400# m1_15000_1400# VSUBS m1_25400_n12200# m1_25400_n2200#
+ m1_25400_400# m1_15000_n8400# m1_25400_n4800# m1_15000_n6000# m1_15000_n1000# m1_25400_n2200#
+ m1_15000_n8400# m1_14840_n13120# m1_15000_n6000# m1_15000_n1000# m1_15000_1400#
+ m1_25400_n9600# m1_15000_n11000# m1_25400_n7200# m1_25400_n7200# m1_25400_n9600#
+ m1_15000_n3400# sky130_fd_pr__res_xhigh_po_5p73_AW8RAB
Xsky130_fd_pr__cap_mim_m3_1_LQXKLG_0 VSUBS m1_15830_n15780# sky130_fd_pr__cap_mim_m3_1_LQXKLG
.ends

.subckt sky130_fd_pr__cap_mim_m3_1_WXTTNJ c1_n2050_n2000# m3_n2150_n2100#
X0 c1_n2050_n2000# m3_n2150_n2100# sky130_fd_pr__cap_mim_m3_1 l=2e+07u w=2e+07u
.ends

.subckt sky130_fd_pr__nfet_01v8_lvt_ZSX9YN a_n210_n643# a_50_n531# a_n50_n557# a_n108_n531#
X0 a_50_n531# a_n50_n557# a_n108_n531# a_n210_n643# sky130_fd_pr__nfet_01v8_lvt ad=1.45e+12p pd=1.058e+07u as=1.45e+12p ps=1.058e+07u w=5e+06u l=500000u
.ends

.subckt sky130_fd_pr__nfet_01v8_lvt_XHV9AV a_50_n281# a_n108_n281# a_n210_n393# a_n50_n307#
X0 a_50_n281# a_n50_n307# a_n108_n281# a_n210_n393# sky130_fd_pr__nfet_01v8_lvt ad=7.25e+11p pd=5.58e+06u as=7.25e+11p ps=5.58e+06u w=2.5e+06u l=500000u
.ends

.subckt sky130_fd_pr__pfet_01v8_TSNZVH a_50_n364# w_n246_n584# a_n108_n364# a_n50_n461#
X0 a_50_n364# a_n50_n461# a_n108_n364# w_n246_n584# sky130_fd_pr__pfet_01v8 ad=1.16e+12p pd=8.58e+06u as=1.16e+12p ps=8.58e+06u w=4e+06u l=500000u
.ends

.subckt sky130_fd_pr__nfet_01v8_Y5UG24 a_n108_n181# a_n50_n207# a_n210_n293# a_50_n181#
X0 a_50_n181# a_n50_n207# a_n108_n181# a_n210_n293# sky130_fd_pr__nfet_01v8 ad=4.35e+11p pd=3.58e+06u as=4.35e+11p ps=3.58e+06u w=1.5e+06u l=500000u
.ends

.subckt inv m1_160_n270# m1_240_n400# li_80_830# VSUBS
Xsky130_fd_pr__pfet_01v8_TSNZVH_0 m1_240_n400# li_80_830# li_80_830# m1_160_n270#
+ sky130_fd_pr__pfet_01v8_TSNZVH
Xsky130_fd_pr__nfet_01v8_Y5UG24_0 VSUBS m1_160_n270# VSUBS m1_240_n400# sky130_fd_pr__nfet_01v8_Y5UG24
.ends

.subckt sample_hold sky130_fd_pr__cap_mim_m3_1_WXTTNJ_0/m3_n2150_n2100# Vcap sky130_fd_pr__nfet_01v8_lvt_ZSX9YN_0/a_50_n531#
+ m1_5220_1840# inv_0/li_80_830# VSUBS
Xsky130_fd_pr__cap_mim_m3_1_WXTTNJ_0 Vcap sky130_fd_pr__cap_mim_m3_1_WXTTNJ_0/m3_n2150_n2100#
+ sky130_fd_pr__cap_mim_m3_1_WXTTNJ
Xsky130_fd_pr__nfet_01v8_lvt_ZSX9YN_0 VSUBS sky130_fd_pr__nfet_01v8_lvt_ZSX9YN_0/a_50_n531#
+ m1_5220_1840# Vcap sky130_fd_pr__nfet_01v8_lvt_ZSX9YN
Xsky130_fd_pr__nfet_01v8_lvt_XHV9AV_0 Vcap Vcap VSUBS m1_5400_600# sky130_fd_pr__nfet_01v8_lvt_XHV9AV
Xinv_0 m1_5220_1840# m1_5400_600# inv_0/li_80_830# VSUBS inv
.ends

.subckt sky130_fd_pr__pfet_01v8_lvt_BKT746 a_287_n764# a_n1451_n764# a_919_n764# w_n1747_n984#
+ a_445_n764# a_1077_n764# a_29_n861# a_603_n764# a_n129_n861# a_187_n861# a_1235_n764#
+ a_n287_n861# a_761_n764# a_819_n861# a_n1077_n861# a_n29_n764# a_345_n861# a_1393_n764#
+ a_n919_n861# a_977_n861# a_n445_n861# a_n187_n764# a_n1235_n861# a_503_n861# a_1551_n764#
+ a_n819_n764# a_1135_n861# a_n603_n861# a_n345_n764# a_n1609_n764# a_661_n861# a_n1393_n861#
+ a_n1135_n764# a_n977_n764# a_1293_n861# a_n761_n861# a_129_n764# a_n503_n764# a_n1293_n764#
+ a_n1551_n861# a_n661_n764# a_1451_n861#
X0 a_n661_n764# a_n761_n861# a_n819_n764# w_n1747_n984# sky130_fd_pr__pfet_01v8_lvt ad=2.32e+12p pd=1.658e+07u as=2.32e+12p ps=1.658e+07u w=8e+06u l=500000u
X1 a_919_n764# a_819_n861# a_761_n764# w_n1747_n984# sky130_fd_pr__pfet_01v8_lvt ad=2.32e+12p pd=1.658e+07u as=2.32e+12p ps=1.658e+07u w=8e+06u l=500000u
X2 a_n187_n764# a_n287_n861# a_n345_n764# w_n1747_n984# sky130_fd_pr__pfet_01v8_lvt ad=2.32e+12p pd=1.658e+07u as=2.32e+12p ps=1.658e+07u w=8e+06u l=500000u
X3 a_761_n764# a_661_n861# a_603_n764# w_n1747_n984# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=2.32e+12p ps=1.658e+07u w=8e+06u l=500000u
X4 a_287_n764# a_187_n861# a_129_n764# w_n1747_n984# sky130_fd_pr__pfet_01v8_lvt ad=2.32e+12p pd=1.658e+07u as=2.32e+12p ps=1.658e+07u w=8e+06u l=500000u
X5 a_n1293_n764# a_n1393_n861# a_n1451_n764# w_n1747_n984# sky130_fd_pr__pfet_01v8_lvt ad=2.32e+12p pd=1.658e+07u as=2.32e+12p ps=1.658e+07u w=8e+06u l=500000u
X6 a_1393_n764# a_1293_n861# a_1235_n764# w_n1747_n984# sky130_fd_pr__pfet_01v8_lvt ad=2.32e+12p pd=1.658e+07u as=2.32e+12p ps=1.658e+07u w=8e+06u l=500000u
X7 a_n345_n764# a_n445_n861# a_n503_n764# w_n1747_n984# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=2.32e+12p ps=1.658e+07u w=8e+06u l=500000u
X8 a_129_n764# a_29_n861# a_n29_n764# w_n1747_n984# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=2.32e+12p ps=1.658e+07u w=8e+06u l=500000u
X9 a_445_n764# a_345_n861# a_287_n764# w_n1747_n984# sky130_fd_pr__pfet_01v8_lvt ad=2.32e+12p pd=1.658e+07u as=0p ps=0u w=8e+06u l=500000u
X10 a_n1451_n764# a_n1551_n861# a_n1609_n764# w_n1747_n984# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=2.32e+12p ps=1.658e+07u w=8e+06u l=500000u
X11 a_1551_n764# a_1451_n861# a_1393_n764# w_n1747_n984# sky130_fd_pr__pfet_01v8_lvt ad=2.32e+12p pd=1.658e+07u as=0p ps=0u w=8e+06u l=500000u
X12 a_n977_n764# a_n1077_n861# a_n1135_n764# w_n1747_n984# sky130_fd_pr__pfet_01v8_lvt ad=2.32e+12p pd=1.658e+07u as=2.32e+12p ps=1.658e+07u w=8e+06u l=500000u
X13 a_n503_n764# a_n603_n861# a_n661_n764# w_n1747_n984# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=8e+06u l=500000u
X14 a_1077_n764# a_977_n861# a_919_n764# w_n1747_n984# sky130_fd_pr__pfet_01v8_lvt ad=2.32e+12p pd=1.658e+07u as=0p ps=0u w=8e+06u l=500000u
X15 a_n29_n764# a_n129_n861# a_n187_n764# w_n1747_n984# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=8e+06u l=500000u
X16 a_603_n764# a_503_n861# a_445_n764# w_n1747_n984# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=8e+06u l=500000u
X17 a_n1135_n764# a_n1235_n861# a_n1293_n764# w_n1747_n984# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=8e+06u l=500000u
X18 a_1235_n764# a_1135_n861# a_1077_n764# w_n1747_n984# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=8e+06u l=500000u
X19 a_n819_n764# a_n919_n861# a_n977_n764# w_n1747_n984# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=8e+06u l=500000u
.ends

.subckt cd_output m1_70_740# sky130_fd_pr__pfet_01v8_lvt_BKT746_0/w_n1747_n984# m1_230_1620#
+ m1_140_70#
Xsky130_fd_pr__pfet_01v8_lvt_BKT746_0 m1_70_740# m1_230_1620# m1_70_740# sky130_fd_pr__pfet_01v8_lvt_BKT746_0/w_n1747_n984#
+ m1_230_1620# m1_230_1620# m1_140_70# m1_70_740# m1_140_70# m1_140_70# m1_70_740#
+ m1_140_70# m1_230_1620# m1_140_70# m1_140_70# m1_70_740# m1_140_70# m1_230_1620#
+ m1_140_70# m1_140_70# m1_140_70# m1_230_1620# m1_140_70# m1_140_70# m1_70_740# m1_230_1620#
+ m1_140_70# m1_140_70# m1_70_740# m1_70_740# m1_140_70# m1_140_70# m1_230_1620# m1_70_740#
+ m1_140_70# m1_140_70# m1_230_1620# m1_230_1620# m1_70_740# m1_140_70# m1_70_740#
+ m1_140_70# sky130_fd_pr__pfet_01v8_lvt_BKT746
.ends

.subckt sky130_fd_pr__pfet_01v8_lvt_D74VRS a_n345_118# a_n661_n1247# a_445_118# a_977_n1344#
+ a_n761_1386# a_n819_1483# a_n345_n2612# a_n819_n2612# a_977_21# a_n977_n1247# a_n345_1483#
+ a_187_21# a_n187_118# a_287_118# a_n187_n2612# a_n1135_1483# a_n977_1483# a_n661_n2612#
+ a_n445_21# a_n819_118# a_n503_1483# a_129_1483# a_919_118# a_n977_n2612# a_n1077_21#
+ a_n661_118# a_761_118# a_29_21# a_345_21# a_29_n2709# a_n661_1483# a_287_1483# a_n603_21#
+ a_29_n1344# a_129_n1247# a_29_1386# a_919_1483# a_603_n1247# a_n129_1386# a_445_1483#
+ a_187_1386# a_n1135_118# a_445_n1247# a_n129_n2709# w_n1273_n2831# a_503_21# a_919_n1247#
+ a_1077_n1247# a_129_n2612# a_1077_1483# a_n603_n2709# a_287_n1247# a_n287_1386#
+ a_n129_n1344# a_819_1386# a_n1077_n2709# a_n977_118# a_1077_118# a_603_n2612# a_n1077_1386#
+ a_603_1483# a_761_n1247# a_n445_n2709# a_503_n2709# a_n29_n1247# a_n919_21# a_n919_n2709#
+ a_345_1386# a_n603_n1344# a_n761_21# a_n129_21# a_129_118# a_445_n2612# a_n919_1386#
+ a_n1077_n1344# a_n287_n2709# a_345_n2709# a_919_n2612# a_819_n2709# a_503_n1344#
+ a_1077_n2612# a_977_1386# a_n445_n1344# a_n445_1386# a_n919_n1344# a_761_1483# a_n1135_n1247#
+ a_n761_n2709# a_287_n2612# a_187_n2709# a_819_21# a_n503_n1247# a_661_21# a_345_n1344#
+ a_n29_118# a_n287_n1344# a_819_n1344# a_503_1386# a_761_n2612# a_n29_1483# a_661_n2709#
+ a_n29_n2612# a_n503_118# a_n761_n1344# a_n345_n1247# a_603_118# a_187_n1344# a_n819_n1247#
+ a_n603_1386# a_n187_1483# a_977_n2709# a_661_n1344# a_n187_n1247# a_661_1386# a_n1135_n2612#
+ a_n287_21# a_n503_n2612#
X0 a_n819_n1247# a_n919_n1344# a_n977_n1247# w_n1273_n2831# sky130_fd_pr__pfet_01v8_lvt ad=1.74e+12p pd=1.258e+07u as=1.74e+12p ps=1.258e+07u w=6e+06u l=500000u
X1 a_n977_n1247# a_n1077_n1344# a_n1135_n1247# w_n1273_n2831# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=1.74e+12p ps=1.258e+07u w=6e+06u l=500000u
X2 a_603_n2612# a_503_n2709# a_445_n2612# w_n1273_n2831# sky130_fd_pr__pfet_01v8_lvt ad=1.74e+12p pd=1.258e+07u as=1.74e+12p ps=1.258e+07u w=6e+06u l=500000u
X3 a_n977_118# a_n1077_21# a_n1135_118# w_n1273_n2831# sky130_fd_pr__pfet_01v8_lvt ad=1.74e+12p pd=1.258e+07u as=1.74e+12p ps=1.258e+07u w=6e+06u l=500000u
X4 a_603_n1247# a_503_n1344# a_445_n1247# w_n1273_n2831# sky130_fd_pr__pfet_01v8_lvt ad=1.74e+12p pd=1.258e+07u as=1.74e+12p ps=1.258e+07u w=6e+06u l=500000u
X5 a_761_n2612# a_661_n2709# a_603_n2612# w_n1273_n2831# sky130_fd_pr__pfet_01v8_lvt ad=1.74e+12p pd=1.258e+07u as=0p ps=0u w=6e+06u l=500000u
X6 a_n819_1483# a_n919_1386# a_n977_1483# w_n1273_n2831# sky130_fd_pr__pfet_01v8_lvt ad=1.74e+12p pd=1.258e+07u as=1.74e+12p ps=1.258e+07u w=6e+06u l=500000u
X7 a_761_n1247# a_661_n1344# a_603_n1247# w_n1273_n2831# sky130_fd_pr__pfet_01v8_lvt ad=1.74e+12p pd=1.258e+07u as=0p ps=0u w=6e+06u l=500000u
X8 a_n661_1483# a_n761_1386# a_n819_1483# w_n1273_n2831# sky130_fd_pr__pfet_01v8_lvt ad=1.74e+12p pd=1.258e+07u as=0p ps=0u w=6e+06u l=500000u
X9 a_919_1483# a_819_1386# a_761_1483# w_n1273_n2831# sky130_fd_pr__pfet_01v8_lvt ad=1.74e+12p pd=1.258e+07u as=1.74e+12p ps=1.258e+07u w=6e+06u l=500000u
X10 a_n187_1483# a_n287_1386# a_n345_1483# w_n1273_n2831# sky130_fd_pr__pfet_01v8_lvt ad=1.74e+12p pd=1.258e+07u as=1.74e+12p ps=1.258e+07u w=6e+06u l=500000u
X11 a_761_1483# a_661_1386# a_603_1483# w_n1273_n2831# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=1.74e+12p ps=1.258e+07u w=6e+06u l=500000u
X12 a_n661_118# a_n761_21# a_n819_118# w_n1273_n2831# sky130_fd_pr__pfet_01v8_lvt ad=1.74e+12p pd=1.258e+07u as=1.74e+12p ps=1.258e+07u w=6e+06u l=500000u
X13 a_n503_n2612# a_n603_n2709# a_n661_n2612# w_n1273_n2831# sky130_fd_pr__pfet_01v8_lvt ad=1.74e+12p pd=1.258e+07u as=1.74e+12p ps=1.258e+07u w=6e+06u l=500000u
X14 a_129_118# a_29_21# a_n29_118# w_n1273_n2831# sky130_fd_pr__pfet_01v8_lvt ad=1.74e+12p pd=1.258e+07u as=1.74e+12p ps=1.258e+07u w=6e+06u l=500000u
X15 a_287_n2612# a_187_n2709# a_129_n2612# w_n1273_n2831# sky130_fd_pr__pfet_01v8_lvt ad=1.74e+12p pd=1.258e+07u as=1.74e+12p ps=1.258e+07u w=6e+06u l=500000u
X16 a_n187_118# a_n287_21# a_n345_118# w_n1273_n2831# sky130_fd_pr__pfet_01v8_lvt ad=1.74e+12p pd=1.258e+07u as=1.74e+12p ps=1.258e+07u w=6e+06u l=500000u
X17 a_n503_n1247# a_n603_n1344# a_n661_n1247# w_n1273_n2831# sky130_fd_pr__pfet_01v8_lvt ad=1.74e+12p pd=1.258e+07u as=1.74e+12p ps=1.258e+07u w=6e+06u l=500000u
X18 a_n661_n2612# a_n761_n2709# a_n819_n2612# w_n1273_n2831# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=1.74e+12p ps=1.258e+07u w=6e+06u l=500000u
X19 a_287_1483# a_187_1386# a_129_1483# w_n1273_n2831# sky130_fd_pr__pfet_01v8_lvt ad=1.74e+12p pd=1.258e+07u as=1.74e+12p ps=1.258e+07u w=6e+06u l=500000u
X20 a_n661_n1247# a_n761_n1344# a_n819_n1247# w_n1273_n2831# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6e+06u l=500000u
X21 a_287_n1247# a_187_n1344# a_129_n1247# w_n1273_n2831# sky130_fd_pr__pfet_01v8_lvt ad=1.74e+12p pd=1.258e+07u as=1.74e+12p ps=1.258e+07u w=6e+06u l=500000u
X22 a_n819_118# a_n919_21# a_n977_118# w_n1273_n2831# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6e+06u l=500000u
X23 a_n345_118# a_n445_21# a_n503_118# w_n1273_n2831# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=1.74e+12p ps=1.258e+07u w=6e+06u l=500000u
X24 a_n503_118# a_n603_21# a_n661_118# w_n1273_n2831# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6e+06u l=500000u
X25 a_n29_n2612# a_n129_n2709# a_n187_n2612# w_n1273_n2831# sky130_fd_pr__pfet_01v8_lvt ad=1.74e+12p pd=1.258e+07u as=1.74e+12p ps=1.258e+07u w=6e+06u l=500000u
X26 a_n345_1483# a_n445_1386# a_n503_1483# w_n1273_n2831# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=1.74e+12p ps=1.258e+07u w=6e+06u l=500000u
X27 a_n29_n1247# a_n129_n1344# a_n187_n1247# w_n1273_n2831# sky130_fd_pr__pfet_01v8_lvt ad=1.74e+12p pd=1.258e+07u as=1.74e+12p ps=1.258e+07u w=6e+06u l=500000u
X28 a_n187_n2612# a_n287_n2709# a_n345_n2612# w_n1273_n2831# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=1.74e+12p ps=1.258e+07u w=6e+06u l=500000u
X29 a_n29_118# a_n129_21# a_n187_118# w_n1273_n2831# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6e+06u l=500000u
X30 a_129_1483# a_29_1386# a_n29_1483# w_n1273_n2831# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=1.74e+12p ps=1.258e+07u w=6e+06u l=500000u
X31 a_n187_n1247# a_n287_n1344# a_n345_n1247# w_n1273_n2831# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=1.74e+12p ps=1.258e+07u w=6e+06u l=500000u
X32 a_445_1483# a_345_1386# a_287_1483# w_n1273_n2831# sky130_fd_pr__pfet_01v8_lvt ad=1.74e+12p pd=1.258e+07u as=0p ps=0u w=6e+06u l=500000u
X33 a_1077_118# a_977_21# a_919_118# w_n1273_n2831# sky130_fd_pr__pfet_01v8_lvt ad=1.74e+12p pd=1.258e+07u as=1.74e+12p ps=1.258e+07u w=6e+06u l=500000u
X34 a_129_n2612# a_29_n2709# a_n29_n2612# w_n1273_n2831# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6e+06u l=500000u
X35 a_n977_1483# a_n1077_1386# a_n1135_1483# w_n1273_n2831# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=1.74e+12p ps=1.258e+07u w=6e+06u l=500000u
X36 a_129_n1247# a_29_n1344# a_n29_n1247# w_n1273_n2831# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6e+06u l=500000u
X37 a_445_n2612# a_345_n2709# a_287_n2612# w_n1273_n2831# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6e+06u l=500000u
X38 a_n503_1483# a_n603_1386# a_n661_1483# w_n1273_n2831# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6e+06u l=500000u
X39 a_1077_1483# a_977_1386# a_919_1483# w_n1273_n2831# sky130_fd_pr__pfet_01v8_lvt ad=1.74e+12p pd=1.258e+07u as=0p ps=0u w=6e+06u l=500000u
X40 a_761_118# a_661_21# a_603_118# w_n1273_n2831# sky130_fd_pr__pfet_01v8_lvt ad=1.74e+12p pd=1.258e+07u as=1.74e+12p ps=1.258e+07u w=6e+06u l=500000u
X41 a_287_118# a_187_21# a_129_118# w_n1273_n2831# sky130_fd_pr__pfet_01v8_lvt ad=1.74e+12p pd=1.258e+07u as=0p ps=0u w=6e+06u l=500000u
X42 a_445_n1247# a_345_n1344# a_287_n1247# w_n1273_n2831# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6e+06u l=500000u
X43 a_919_n2612# a_819_n2709# a_761_n2612# w_n1273_n2831# sky130_fd_pr__pfet_01v8_lvt ad=1.74e+12p pd=1.258e+07u as=0p ps=0u w=6e+06u l=500000u
X44 a_n29_1483# a_n129_1386# a_n187_1483# w_n1273_n2831# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6e+06u l=500000u
X45 a_603_1483# a_503_1386# a_445_1483# w_n1273_n2831# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6e+06u l=500000u
X46 a_445_118# a_345_21# a_287_118# w_n1273_n2831# sky130_fd_pr__pfet_01v8_lvt ad=1.74e+12p pd=1.258e+07u as=0p ps=0u w=6e+06u l=500000u
X47 a_919_118# a_819_21# a_761_118# w_n1273_n2831# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6e+06u l=500000u
X48 a_919_n1247# a_819_n1344# a_761_n1247# w_n1273_n2831# sky130_fd_pr__pfet_01v8_lvt ad=1.74e+12p pd=1.258e+07u as=0p ps=0u w=6e+06u l=500000u
X49 a_1077_n2612# a_977_n2709# a_919_n2612# w_n1273_n2831# sky130_fd_pr__pfet_01v8_lvt ad=1.74e+12p pd=1.258e+07u as=0p ps=0u w=6e+06u l=500000u
X50 a_1077_n1247# a_977_n1344# a_919_n1247# w_n1273_n2831# sky130_fd_pr__pfet_01v8_lvt ad=1.74e+12p pd=1.258e+07u as=0p ps=0u w=6e+06u l=500000u
X51 a_603_118# a_503_21# a_445_118# w_n1273_n2831# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6e+06u l=500000u
X52 a_n345_n2612# a_n445_n2709# a_n503_n2612# w_n1273_n2831# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6e+06u l=500000u
X53 a_n345_n1247# a_n445_n1344# a_n503_n1247# w_n1273_n2831# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6e+06u l=500000u
X54 a_n819_n2612# a_n919_n2709# a_n977_n2612# w_n1273_n2831# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=1.74e+12p ps=1.258e+07u w=6e+06u l=500000u
X55 a_n977_n2612# a_n1077_n2709# a_n1135_n2612# w_n1273_n2831# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=1.74e+12p ps=1.258e+07u w=6e+06u l=500000u
.ends

.subckt XM_cs li_876_5462# m1_52_164# m1_147_79#
Xsky130_fd_pr__pfet_01v8_lvt_D74VRS_0 li_876_5462# li_876_5462# m1_52_164# m1_147_79#
+ m1_147_79# m1_52_164# li_876_5462# m1_52_164# m1_147_79# li_876_5462# li_876_5462#
+ m1_147_79# m1_52_164# li_876_5462# m1_52_164# m1_52_164# li_876_5462# li_876_5462#
+ m1_147_79# m1_52_164# m1_52_164# m1_52_164# li_876_5462# li_876_5462# m1_147_79#
+ li_876_5462# m1_52_164# m1_147_79# m1_147_79# m1_147_79# li_876_5462# li_876_5462#
+ m1_147_79# m1_147_79# m1_52_164# m1_147_79# li_876_5462# li_876_5462# m1_147_79#
+ m1_52_164# m1_147_79# m1_52_164# m1_52_164# m1_147_79# li_876_5462# m1_147_79# li_876_5462#
+ m1_52_164# m1_52_164# m1_52_164# m1_147_79# li_876_5462# m1_147_79# m1_147_79# m1_147_79#
+ m1_147_79# li_876_5462# m1_52_164# li_876_5462# m1_147_79# li_876_5462# m1_52_164#
+ m1_147_79# m1_147_79# li_876_5462# m1_147_79# m1_147_79# m1_147_79# m1_147_79# m1_147_79#
+ m1_147_79# m1_52_164# m1_52_164# m1_147_79# m1_147_79# m1_147_79# m1_147_79# li_876_5462#
+ m1_147_79# m1_147_79# m1_52_164# m1_147_79# m1_147_79# m1_147_79# m1_147_79# m1_52_164#
+ m1_52_164# m1_147_79# li_876_5462# m1_147_79# m1_147_79# m1_52_164# m1_147_79# m1_147_79#
+ li_876_5462# m1_147_79# m1_147_79# m1_147_79# m1_52_164# li_876_5462# m1_147_79#
+ li_876_5462# m1_52_164# m1_147_79# li_876_5462# li_876_5462# m1_147_79# m1_52_164#
+ m1_147_79# m1_52_164# m1_147_79# m1_147_79# m1_52_164# m1_147_79# m1_52_164# m1_147_79#
+ m1_52_164# sky130_fd_pr__pfet_01v8_lvt_D74VRS
.ends

.subckt sky130_fd_pr__nfet_01v8_lvt_E96B6C a_29_n507# a_n287_n419# a_n229_n507# a_287_n507#
+ a_229_n419# a_n545_n419# a_n487_n507# a_n29_n419# a_487_n419# VSUBS
X0 a_487_n419# a_287_n507# a_229_n419# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=1.305e+12p pd=9.58e+06u as=1.305e+12p ps=9.58e+06u w=4.5e+06u l=1e+06u
X1 a_n29_n419# a_n229_n507# a_n287_n419# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=1.305e+12p pd=9.58e+06u as=1.305e+12p ps=9.58e+06u w=4.5e+06u l=1e+06u
X2 a_229_n419# a_29_n507# a_n29_n419# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4.5e+06u l=1e+06u
X3 a_n287_n419# a_n487_n507# a_n545_n419# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=1.305e+12p ps=9.58e+06u w=4.5e+06u l=1e+06u
.ends

.subckt sky130_fd_pr__nfet_01v8_lvt_A5VCMN a_229_n481# a_29_n507# a_n545_n481# a_n229_n507#
+ a_287_n507# a_n29_n481# a_487_n481# a_n487_n507# a_n287_n481# VSUBS
X0 a_487_n481# a_287_n507# a_229_n481# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=1.305e+12p pd=9.58e+06u as=1.305e+12p ps=9.58e+06u w=4.5e+06u l=1e+06u
X1 a_229_n481# a_29_n507# a_n29_n481# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=1.305e+12p ps=9.58e+06u w=4.5e+06u l=1e+06u
X2 a_n29_n481# a_n229_n507# a_n287_n481# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=1.305e+12p ps=9.58e+06u w=4.5e+06u l=1e+06u
X3 a_n287_n481# a_n487_n507# a_n545_n481# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=1.305e+12p ps=9.58e+06u w=4.5e+06u l=1e+06u
.ends

.subckt XM_diffpair m1_160_200# sky130_fd_pr__nfet_01v8_lvt_E96B6C_0/VSUBS m1_30_1280#
+ m1_30_n1060# m1_280_n670# m1_551_360#
Xsky130_fd_pr__nfet_01v8_lvt_E96B6C_0 m1_551_360# m1_280_n670# m1_551_360# m1_160_200#
+ m1_280_n670# m1_30_1280# m1_160_200# m1_30_n1060# m1_30_1280# sky130_fd_pr__nfet_01v8_lvt_E96B6C_0/VSUBS
+ sky130_fd_pr__nfet_01v8_lvt_E96B6C
Xsky130_fd_pr__nfet_01v8_lvt_A5VCMN_0 m1_280_n670# m1_160_200# m1_30_n1060# m1_160_200#
+ m1_551_360# m1_30_1280# m1_30_n1060# m1_551_360# m1_280_n670# sky130_fd_pr__nfet_01v8_lvt_E96B6C_0/VSUBS
+ sky130_fd_pr__nfet_01v8_lvt_A5VCMN
.ends

.subckt sky130_fd_pr__cap_mim_m3_1_EN3Q86 c1_n1650_n2140# m3_n1750_n2240#
X0 c1_n1650_n2140# m3_n1750_n2240# sky130_fd_pr__cap_mim_m3_1 l=2.14e+07u w=1.6e+07u
.ends

.subckt sky130_fd_pr__res_high_po_2p85_7J2RPB a_n285_n1642# a_n415_n1772# a_n285_1210#
X0 a_n285_n1642# a_n285_1210# a_n415_n1772# sky130_fd_pr__res_high_po_2p85 l=1.21e+07u
.ends

.subckt sky130_fd_pr__nfet_01v8_lvt_USQY94 a_n1174_n1403# a_658_109# a_n716_n1403#
+ a_200_109# a_n1116_21# a_1116_865# a_n258_n1403# a_n200_n1491# a_716_n1491# a_n1174_n647#
+ a_n200_21# a_n658_n1491# a_n200_n735# a_n258_865# a_1116_109# a_200_n647# a_258_21#
+ a_n658_21# a_1116_n1403# a_258_n1491# a_258_777# a_n1276_n1577# a_n1116_n735# a_n258_109#
+ a_n716_n647# a_n1174_865# a_n658_777# a_n200_777# a_n258_n647# a_n716_865# a_n658_n735#
+ a_200_n1403# a_1116_n647# a_n1174_109# a_716_21# a_658_n1403# a_716_n735# a_658_865#
+ a_716_777# a_658_n647# a_258_n735# a_200_865# a_n1116_n1491# a_n716_109# a_n1116_777#
X0 a_658_n1403# a_258_n1491# a_200_n1403# a_n1276_n1577# sky130_fd_pr__nfet_01v8_lvt ad=8.7e+11p pd=6.58e+06u as=8.7e+11p ps=6.58e+06u w=3e+06u l=2e+06u
X1 a_n716_n1403# a_n1116_n1491# a_n1174_n1403# a_n1276_n1577# sky130_fd_pr__nfet_01v8_lvt ad=8.7e+11p pd=6.58e+06u as=8.7e+11p ps=6.58e+06u w=3e+06u l=2e+06u
X2 a_658_109# a_258_21# a_200_109# a_n1276_n1577# sky130_fd_pr__nfet_01v8_lvt ad=8.7e+11p pd=6.58e+06u as=8.7e+11p ps=6.58e+06u w=3e+06u l=2e+06u
X3 a_1116_n647# a_716_n735# a_658_n647# a_n1276_n1577# sky130_fd_pr__nfet_01v8_lvt ad=8.7e+11p pd=6.58e+06u as=8.7e+11p ps=6.58e+06u w=3e+06u l=2e+06u
X4 a_1116_n1403# a_716_n1491# a_658_n1403# a_n1276_n1577# sky130_fd_pr__nfet_01v8_lvt ad=8.7e+11p pd=6.58e+06u as=0p ps=0u w=3e+06u l=2e+06u
X5 a_200_865# a_n200_777# a_n258_865# a_n1276_n1577# sky130_fd_pr__nfet_01v8_lvt ad=8.7e+11p pd=6.58e+06u as=8.7e+11p ps=6.58e+06u w=3e+06u l=2e+06u
X6 a_1116_109# a_716_21# a_658_109# a_n1276_n1577# sky130_fd_pr__nfet_01v8_lvt ad=8.7e+11p pd=6.58e+06u as=0p ps=0u w=3e+06u l=2e+06u
X7 a_200_n647# a_n200_n735# a_n258_n647# a_n1276_n1577# sky130_fd_pr__nfet_01v8_lvt ad=8.7e+11p pd=6.58e+06u as=8.7e+11p ps=6.58e+06u w=3e+06u l=2e+06u
X8 a_n716_n647# a_n1116_n735# a_n1174_n647# a_n1276_n1577# sky130_fd_pr__nfet_01v8_lvt ad=8.7e+11p pd=6.58e+06u as=8.7e+11p ps=6.58e+06u w=3e+06u l=2e+06u
X9 a_n258_865# a_n658_777# a_n716_865# a_n1276_n1577# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=8.7e+11p ps=6.58e+06u w=3e+06u l=2e+06u
X10 a_n716_865# a_n1116_777# a_n1174_865# a_n1276_n1577# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=8.7e+11p ps=6.58e+06u w=3e+06u l=2e+06u
X11 a_658_n647# a_258_n735# a_200_n647# a_n1276_n1577# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=2e+06u
X12 a_200_109# a_n200_21# a_n258_109# a_n1276_n1577# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=8.7e+11p ps=6.58e+06u w=3e+06u l=2e+06u
X13 a_658_865# a_258_777# a_200_865# a_n1276_n1577# sky130_fd_pr__nfet_01v8_lvt ad=8.7e+11p pd=6.58e+06u as=0p ps=0u w=3e+06u l=2e+06u
X14 a_n258_109# a_n658_21# a_n716_109# a_n1276_n1577# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=8.7e+11p ps=6.58e+06u w=3e+06u l=2e+06u
X15 a_n258_n647# a_n658_n735# a_n716_n647# a_n1276_n1577# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=2e+06u
X16 a_200_n1403# a_n200_n1491# a_n258_n1403# a_n1276_n1577# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=8.7e+11p ps=6.58e+06u w=3e+06u l=2e+06u
X17 a_1116_865# a_716_777# a_658_865# a_n1276_n1577# sky130_fd_pr__nfet_01v8_lvt ad=8.7e+11p pd=6.58e+06u as=0p ps=0u w=3e+06u l=2e+06u
X18 a_n716_109# a_n1116_21# a_n1174_109# a_n1276_n1577# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=8.7e+11p ps=6.58e+06u w=3e+06u l=2e+06u
X19 a_n258_n1403# a_n658_n1491# a_n716_n1403# a_n1276_n1577# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=2e+06u
.ends

.subckt XM_actload2 m1_985_79# m1_522_658# m1_522_1414# m1_62_1668# m1_522_2926# m1_520_2170#
+ VSUBS
Xsky130_fd_pr__nfet_01v8_lvt_USQY94_0 m1_62_1668# m1_62_1668# m1_522_658# m1_520_2170#
+ m1_985_79# m1_522_2926# m1_62_1668# m1_985_79# m1_985_79# m1_62_1668# m1_985_79#
+ m1_985_79# m1_985_79# m1_62_1668# m1_520_2170# m1_522_1414# m1_985_79# m1_985_79#
+ m1_522_658# m1_985_79# m1_985_79# VSUBS m1_985_79# m1_62_1668# m1_522_1414# m1_62_1668#
+ m1_985_79# m1_985_79# m1_62_1668# m1_522_2926# m1_985_79# m1_522_658# m1_522_1414#
+ m1_62_1668# m1_985_79# m1_62_1668# m1_985_79# m1_62_1668# m1_985_79# m1_62_1668#
+ m1_985_79# m1_522_2926# m1_985_79# m1_520_2170# m1_985_79# sky130_fd_pr__nfet_01v8_lvt_USQY94
.ends

.subckt sky130_fd_pr__nfet_01v8_lvt_7MFZYU a_n429_299# a_29_299# a_n487_n725# a_429_387#
+ a_429_n1281# a_n29_n725# a_n487_943# a_n429_n813# a_429_n725# a_n487_n169# a_29_n813#
+ a_n29_943# a_n589_n1455# a_29_n1369# a_n29_n1281# a_n29_n169# a_n487_387# a_n429_n257#
+ a_29_855# a_n429_855# a_n429_n1369# a_429_n169# a_n487_n1281# a_29_n257# a_n29_387#
+ a_429_943#
X0 a_429_n169# a_29_n257# a_n29_n169# a_n589_n1455# sky130_fd_pr__nfet_01v8_lvt ad=5.8e+11p pd=4.58e+06u as=5.8e+11p ps=4.58e+06u w=2e+06u l=2e+06u
X1 a_429_n725# a_29_n813# a_n29_n725# a_n589_n1455# sky130_fd_pr__nfet_01v8_lvt ad=5.8e+11p pd=4.58e+06u as=5.8e+11p ps=4.58e+06u w=2e+06u l=2e+06u
X2 a_n29_n1281# a_n429_n1369# a_n487_n1281# a_n589_n1455# sky130_fd_pr__nfet_01v8_lvt ad=5.8e+11p pd=4.58e+06u as=5.8e+11p ps=4.58e+06u w=2e+06u l=2e+06u
X3 a_429_387# a_29_299# a_n29_387# a_n589_n1455# sky130_fd_pr__nfet_01v8_lvt ad=5.8e+11p pd=4.58e+06u as=5.8e+11p ps=4.58e+06u w=2e+06u l=2e+06u
X4 a_429_943# a_29_855# a_n29_943# a_n589_n1455# sky130_fd_pr__nfet_01v8_lvt ad=5.8e+11p pd=4.58e+06u as=5.8e+11p ps=4.58e+06u w=2e+06u l=2e+06u
X5 a_429_n1281# a_29_n1369# a_n29_n1281# a_n589_n1455# sky130_fd_pr__nfet_01v8_lvt ad=5.8e+11p pd=4.58e+06u as=0p ps=0u w=2e+06u l=2e+06u
X6 a_n29_n169# a_n429_n257# a_n487_n169# a_n589_n1455# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=5.8e+11p ps=4.58e+06u w=2e+06u l=2e+06u
X7 a_n29_n725# a_n429_n813# a_n487_n725# a_n589_n1455# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=5.8e+11p ps=4.58e+06u w=2e+06u l=2e+06u
X8 a_n29_943# a_n429_855# a_n487_943# a_n589_n1455# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=5.8e+11p ps=4.58e+06u w=2e+06u l=2e+06u
X9 a_n29_387# a_n429_299# a_n487_387# a_n589_n1455# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=5.8e+11p ps=4.58e+06u w=2e+06u l=2e+06u
.ends

.subckt XM_tail m1_530_330# m1_780_80# VSUBS
Xsky130_fd_pr__nfet_01v8_lvt_7MFZYU_0 m1_780_80# m1_780_80# VSUBS VSUBS VSUBS m1_530_330#
+ VSUBS m1_780_80# VSUBS VSUBS m1_780_80# m1_530_330# VSUBS m1_780_80# m1_530_330#
+ m1_530_330# VSUBS m1_780_80# m1_780_80# m1_780_80# m1_780_80# VSUBS VSUBS m1_780_80#
+ m1_530_330# VSUBS sky130_fd_pr__nfet_01v8_lvt_7MFZYU
.ends

.subckt sky130_fd_pr__pfet_01v8_lvt_MBDTEX a_745_n236# a_545_n262# a_1777_n236# a_1577_n262#
+ a_229_n236# a_n1577_n236# a_2035_n236# a_n1777_n262# a_29_n262# w_n2129_n298# a_n545_n236#
+ a_n745_n262# a_1003_n236# a_803_n262# a_n2035_n262# a_1835_n262# a_n29_n236# a_n229_n262#
+ a_487_n236# a_287_n262# a_n1003_n262# a_n1835_n236# a_n803_n236# a_1519_n236# a_n2093_n236#
+ a_1319_n262# a_1261_n236# a_1061_n262# a_n1319_n236# a_n287_n236# a_n1061_n236#
+ a_n1519_n262# a_n487_n262# a_n1261_n262#
X0 a_n1061_n236# a_n1261_n262# a_n1319_n236# w_n2129_n298# sky130_fd_pr__pfet_01v8_lvt ad=5.8e+11p pd=4.58e+06u as=5.8e+11p ps=4.58e+06u w=2e+06u l=1e+06u
X1 a_745_n236# a_545_n262# a_487_n236# w_n2129_n298# sky130_fd_pr__pfet_01v8_lvt ad=5.8e+11p pd=4.58e+06u as=5.8e+11p ps=4.58e+06u w=2e+06u l=1e+06u
X2 a_1003_n236# a_803_n262# a_745_n236# w_n2129_n298# sky130_fd_pr__pfet_01v8_lvt ad=5.8e+11p pd=4.58e+06u as=0p ps=0u w=2e+06u l=1e+06u
X3 a_487_n236# a_287_n262# a_229_n236# w_n2129_n298# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=5.8e+11p ps=4.58e+06u w=2e+06u l=1e+06u
X4 a_2035_n236# a_1835_n262# a_1777_n236# w_n2129_n298# sky130_fd_pr__pfet_01v8_lvt ad=5.8e+11p pd=4.58e+06u as=5.8e+11p ps=4.58e+06u w=2e+06u l=1e+06u
X5 a_1777_n236# a_1577_n262# a_1519_n236# w_n2129_n298# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=5.8e+11p ps=4.58e+06u w=2e+06u l=1e+06u
X6 a_1261_n236# a_1061_n262# a_1003_n236# w_n2129_n298# sky130_fd_pr__pfet_01v8_lvt ad=5.8e+11p pd=4.58e+06u as=0p ps=0u w=2e+06u l=1e+06u
X7 a_n1835_n236# a_n2035_n262# a_n2093_n236# w_n2129_n298# sky130_fd_pr__pfet_01v8_lvt ad=5.8e+11p pd=4.58e+06u as=5.8e+11p ps=4.58e+06u w=2e+06u l=1e+06u
X8 a_n29_n236# a_n229_n262# a_n287_n236# w_n2129_n298# sky130_fd_pr__pfet_01v8_lvt ad=5.8e+11p pd=4.58e+06u as=5.8e+11p ps=4.58e+06u w=2e+06u l=1e+06u
X9 a_229_n236# a_29_n262# a_n29_n236# w_n2129_n298# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X10 a_n1319_n236# a_n1519_n262# a_n1577_n236# w_n2129_n298# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=5.8e+11p ps=4.58e+06u w=2e+06u l=1e+06u
X11 a_n545_n236# a_n745_n262# a_n803_n236# w_n2129_n298# sky130_fd_pr__pfet_01v8_lvt ad=5.8e+11p pd=4.58e+06u as=5.8e+11p ps=4.58e+06u w=2e+06u l=1e+06u
X12 a_n803_n236# a_n1003_n262# a_n1061_n236# w_n2129_n298# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X13 a_n287_n236# a_n487_n262# a_n545_n236# w_n2129_n298# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X14 a_n1577_n236# a_n1777_n262# a_n1835_n236# w_n2129_n298# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X15 a_1519_n236# a_1319_n262# a_1261_n236# w_n2129_n298# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
.ends

.subckt sky130_fd_pr__pfet_01v8_lvt_B64SAM a_545_n261# a_1777_n164# a_1577_n261# a_229_n164#
+ a_n1577_n164# a_2035_n164# a_n545_n164# a_29_n261# a_n1777_n261# a_n745_n261# a_1003_n164#
+ a_803_n261# a_n2035_n261# a_n29_n164# a_487_n164# a_1835_n261# a_n229_n261# w_n2129_n264#
+ a_n1835_n164# a_287_n261# a_n1003_n261# a_n803_n164# a_1519_n164# a_n2093_n164#
+ a_1261_n164# a_1319_n261# a_n1319_n164# a_1061_n261# a_n287_n164# a_n1061_n164#
+ a_n1519_n261# a_745_n164# a_n487_n261# a_n1261_n261#
X0 a_n29_n164# a_n229_n261# a_n287_n164# w_n2129_n264# sky130_fd_pr__pfet_01v8_lvt ad=5.8e+11p pd=4.58e+06u as=5.8e+11p ps=4.58e+06u w=2e+06u l=1e+06u
X1 a_229_n164# a_29_n261# a_n29_n164# w_n2129_n264# sky130_fd_pr__pfet_01v8_lvt ad=5.8e+11p pd=4.58e+06u as=0p ps=0u w=2e+06u l=1e+06u
X2 a_n1319_n164# a_n1519_n261# a_n1577_n164# w_n2129_n264# sky130_fd_pr__pfet_01v8_lvt ad=5.8e+11p pd=4.58e+06u as=5.8e+11p ps=4.58e+06u w=2e+06u l=1e+06u
X3 a_n545_n164# a_n745_n261# a_n803_n164# w_n2129_n264# sky130_fd_pr__pfet_01v8_lvt ad=5.8e+11p pd=4.58e+06u as=5.8e+11p ps=4.58e+06u w=2e+06u l=1e+06u
X4 a_n287_n164# a_n487_n261# a_n545_n164# w_n2129_n264# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X5 a_n803_n164# a_n1003_n261# a_n1061_n164# w_n2129_n264# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=5.8e+11p ps=4.58e+06u w=2e+06u l=1e+06u
X6 a_n1577_n164# a_n1777_n261# a_n1835_n164# w_n2129_n264# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=5.8e+11p ps=4.58e+06u w=2e+06u l=1e+06u
X7 a_1519_n164# a_1319_n261# a_1261_n164# w_n2129_n264# sky130_fd_pr__pfet_01v8_lvt ad=5.8e+11p pd=4.58e+06u as=5.8e+11p ps=4.58e+06u w=2e+06u l=1e+06u
X8 a_n1061_n164# a_n1261_n261# a_n1319_n164# w_n2129_n264# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X9 a_1003_n164# a_803_n261# a_745_n164# w_n2129_n264# sky130_fd_pr__pfet_01v8_lvt ad=5.8e+11p pd=4.58e+06u as=5.8e+11p ps=4.58e+06u w=2e+06u l=1e+06u
X10 a_745_n164# a_545_n261# a_487_n164# w_n2129_n264# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=5.8e+11p ps=4.58e+06u w=2e+06u l=1e+06u
X11 a_487_n164# a_287_n261# a_229_n164# w_n2129_n264# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X12 a_1777_n164# a_1577_n261# a_1519_n164# w_n2129_n264# sky130_fd_pr__pfet_01v8_lvt ad=5.8e+11p pd=4.58e+06u as=0p ps=0u w=2e+06u l=1e+06u
X13 a_2035_n164# a_1835_n261# a_1777_n164# w_n2129_n264# sky130_fd_pr__pfet_01v8_lvt ad=5.8e+11p pd=4.58e+06u as=0p ps=0u w=2e+06u l=1e+06u
X14 a_1261_n164# a_1061_n261# a_1003_n164# w_n2129_n264# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X15 a_n1835_n164# a_n2035_n261# a_n2093_n164# w_n2129_n264# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=5.8e+11p ps=4.58e+06u w=2e+06u l=1e+06u
.ends

.subckt XM_ppair w_n220_n1060# m1_240_n480# m1_70_n360#
Xsky130_fd_pr__pfet_01v8_lvt_MBDTEX_0 m1_70_n360# m1_70_n360# m1_240_n480# m1_70_n360#
+ m1_240_n480# w_n220_n1060# w_n220_n1060# m1_70_n360# m1_70_n360# w_n220_n1060# w_n220_n1060#
+ m1_70_n360# w_n220_n1060# m1_70_n360# m1_70_n360# m1_70_n360# w_n220_n1060# m1_70_n360#
+ w_n220_n1060# m1_70_n360# m1_70_n360# m1_240_n480# m1_70_n360# w_n220_n1060# w_n220_n1060#
+ m1_70_n360# m1_70_n360# m1_70_n360# m1_70_n360# m1_240_n480# w_n220_n1060# m1_70_n360#
+ m1_70_n360# m1_70_n360# sky130_fd_pr__pfet_01v8_lvt_MBDTEX
Xsky130_fd_pr__pfet_01v8_lvt_B64SAM_0 m1_70_n360# m1_70_n360# m1_70_n360# m1_70_n360#
+ w_n220_n1060# w_n220_n1060# w_n220_n1060# m1_70_n360# m1_70_n360# m1_70_n360# w_n220_n1060#
+ m1_70_n360# m1_70_n360# w_n220_n1060# w_n220_n1060# m1_70_n360# m1_70_n360# w_n220_n1060#
+ m1_70_n360# m1_70_n360# m1_70_n360# m1_240_n480# w_n220_n1060# w_n220_n1060# m1_240_n480#
+ m1_70_n360# m1_240_n480# m1_70_n360# m1_70_n360# w_n220_n1060# m1_70_n360# m1_240_n480#
+ m1_70_n360# m1_70_n360# sky130_fd_pr__pfet_01v8_lvt_B64SAM
.ends

.subckt opamp_realcomp3_usefinger in_n in_p bias_0p7 out vdd vss
XXM_cs_0 vdd out first_stage_out XM_cs
XXM_diffpair_0 in_p vss first_stage_out ppair_gate m2_n4080_2260# in_n XM_diffpair
Xsky130_fd_pr__cap_mim_m3_1_EN3Q86_0 first_stage_out m1_6290_1100# sky130_fd_pr__cap_mim_m3_1_EN3Q86
Xsky130_fd_pr__res_high_po_2p85_7J2RPB_0 out vss m1_6290_1100# sky130_fd_pr__res_high_po_2p85_7J2RPB
XXM_actload2_0 bias_0p7 out out vss out out vss XM_actload2
XXM_tail_0 m2_n4080_2260# bias_0p7 vss XM_tail
XXM_ppair_0 vdd first_stage_out ppair_gate XM_ppair
.ends

.subckt sky130_fd_pr__nfet_01v8_lvt_J9QE6F a_n2548_n69# a_716_n157# a_2490_n69# a_258_n157#
+ a_n258_n69# a_n2490_n157# a_2032_n69# a_n2032_n157# a_n2650_n243# a_n1174_n69# a_n716_n69#
+ a_2090_n157# a_n200_n157# a_658_n69# a_n1574_n157# a_n2090_n69# a_200_n69# a_n1116_n157#
+ a_n1632_n69# a_1574_n69# a_1632_n157# a_1174_n157# a_1116_n69# a_n658_n157#
X0 a_658_n69# a_258_n157# a_200_n69# a_n2650_n243# sky130_fd_pr__nfet_01v8_lvt ad=2.9e+11p pd=2.58e+06u as=2.9e+11p ps=2.58e+06u w=1e+06u l=2e+06u
X1 a_2490_n69# a_2090_n157# a_2032_n69# a_n2650_n243# sky130_fd_pr__nfet_01v8_lvt ad=2.9e+11p pd=2.58e+06u as=2.9e+11p ps=2.58e+06u w=1e+06u l=2e+06u
X2 a_1574_n69# a_1174_n157# a_1116_n69# a_n2650_n243# sky130_fd_pr__nfet_01v8_lvt ad=2.9e+11p pd=2.58e+06u as=2.9e+11p ps=2.58e+06u w=1e+06u l=2e+06u
X3 a_1116_n69# a_716_n157# a_658_n69# a_n2650_n243# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X4 a_2032_n69# a_1632_n157# a_1574_n69# a_n2650_n243# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X5 a_200_n69# a_n200_n157# a_n258_n69# a_n2650_n243# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=2.9e+11p ps=2.58e+06u w=1e+06u l=2e+06u
X6 a_n2090_n69# a_n2490_n157# a_n2548_n69# a_n2650_n243# sky130_fd_pr__nfet_01v8_lvt ad=2.9e+11p pd=2.58e+06u as=2.9e+11p ps=2.58e+06u w=1e+06u l=2e+06u
X7 a_n1632_n69# a_n2032_n157# a_n2090_n69# a_n2650_n243# sky130_fd_pr__nfet_01v8_lvt ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=2e+06u
X8 a_n1174_n69# a_n1574_n157# a_n1632_n69# a_n2650_n243# sky130_fd_pr__nfet_01v8_lvt ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=2e+06u
X9 a_n258_n69# a_n658_n157# a_n716_n69# a_n2650_n243# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=2.9e+11p ps=2.58e+06u w=1e+06u l=2e+06u
X10 a_n716_n69# a_n1116_n157# a_n1174_n69# a_n2650_n243# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
.ends

.subckt sky130_fd_pr__nfet_01v8_lvt_M93XMJ a_716_n157# a_258_n157# a_n2490_n157# a_2490_n131#
+ a_n1632_n131# a_n2032_n157# a_n1174_n131# a_n2548_n131# a_2032_n131# a_n2650_n243#
+ a_200_n131# a_2090_n157# a_n200_n157# a_n716_n131# a_n1574_n157# a_n258_n131# a_1574_n131#
+ a_n1116_n157# a_1116_n131# a_n2090_n131# a_1632_n157# a_658_n131# a_1174_n157# a_n658_n157#
X0 a_200_n131# a_n200_n157# a_n258_n131# a_n2650_n243# sky130_fd_pr__nfet_01v8_lvt ad=2.9e+11p pd=2.58e+06u as=2.9e+11p ps=2.58e+06u w=1e+06u l=2e+06u
X1 a_2032_n131# a_1632_n157# a_1574_n131# a_n2650_n243# sky130_fd_pr__nfet_01v8_lvt ad=2.9e+11p pd=2.58e+06u as=2.9e+11p ps=2.58e+06u w=1e+06u l=2e+06u
X2 a_n716_n131# a_n1116_n157# a_n1174_n131# a_n2650_n243# sky130_fd_pr__nfet_01v8_lvt ad=2.9e+11p pd=2.58e+06u as=2.9e+11p ps=2.58e+06u w=1e+06u l=2e+06u
X3 a_2490_n131# a_2090_n157# a_2032_n131# a_n2650_n243# sky130_fd_pr__nfet_01v8_lvt ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=2e+06u
X4 a_n2090_n131# a_n2490_n157# a_n2548_n131# a_n2650_n243# sky130_fd_pr__nfet_01v8_lvt ad=2.9e+11p pd=2.58e+06u as=2.9e+11p ps=2.58e+06u w=1e+06u l=2e+06u
X5 a_658_n131# a_258_n157# a_200_n131# a_n2650_n243# sky130_fd_pr__nfet_01v8_lvt ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=2e+06u
X6 a_n258_n131# a_n658_n157# a_n716_n131# a_n2650_n243# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X7 a_1574_n131# a_1174_n157# a_1116_n131# a_n2650_n243# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=2.9e+11p ps=2.58e+06u w=1e+06u l=2e+06u
X8 a_n1632_n131# a_n2032_n157# a_n2090_n131# a_n2650_n243# sky130_fd_pr__nfet_01v8_lvt ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=2e+06u
X9 a_n1174_n131# a_n1574_n157# a_n1632_n131# a_n2650_n243# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X10 a_1116_n131# a_716_n157# a_658_n131# a_n2650_n243# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
.ends

.subckt cd_current m1_1080_160# m1_1080_870# m1_1070_700# VSUBS
Xsky130_fd_pr__nfet_01v8_lvt_J9QE6F_1 VSUBS m1_1080_160# VSUBS m1_1080_160# m1_640_380#
+ VSUBS VSUBS m1_1080_160# VSUBS m1_640_380# VSUBS VSUBS m1_1080_160# m1_640_380#
+ m1_1080_160# m1_640_380# VSUBS m1_1080_160# VSUBS m1_640_380# m1_1080_160# m1_1080_160#
+ VSUBS m1_1080_160# sky130_fd_pr__nfet_01v8_lvt_J9QE6F
Xsky130_fd_pr__nfet_01v8_lvt_M93XMJ_0 m1_1080_870# m1_1080_870# VSUBS VSUBS m1_1070_700#
+ m1_1080_870# m1_640_380# VSUBS m1_1070_700# VSUBS m1_1070_700# VSUBS m1_1080_870#
+ m1_1070_700# m1_1080_870# m1_640_380# m1_640_380# m1_1080_870# m1_1070_700# m1_640_380#
+ m1_1080_870# m1_640_380# m1_1080_870# m1_1080_870# sky130_fd_pr__nfet_01v8_lvt_M93XMJ
.ends

.subckt sky130_fd_pr__pfet_01v8_lvt_QH9SH3 a_n2548_118# a_2490_118# a_n258_118# a_1116_n3318#
+ a_n1116_21# w_n2686_n3537# a_2032_118# a_1574_n3318# a_2032_n3318# a_n1116_n3415#
+ a_n200_21# a_n2032_21# a_n1174_118# a_n1574_n3415# a_2490_n3318# a_200_n3318# a_n1632_n3318#
+ a_1632_n3415# a_n716_118# a_n2032_n3415# a_258_21# a_n658_21# a_658_n3318# a_n1574_21#
+ a_n2548_n3318# a_n2490_n3415# a_658_118# a_1174_21# a_n2090_118# a_n1174_n3318#
+ a_1174_n3415# a_200_118# a_n200_n3415# a_716_n3415# a_n658_n3415# a_n1632_118# a_n2490_21#
+ a_2090_21# a_n716_n3318# a_n2090_n3318# a_2090_n3415# a_1574_118# a_716_21# a_258_n3415#
+ a_1632_21# a_1116_118# a_n258_n3318#
X0 a_n1632_118# a_n2032_21# a_n2090_118# w_n2686_n3537# sky130_fd_pr__pfet_01v8_lvt ad=4.64e+12p pd=3.258e+07u as=4.64e+12p ps=3.258e+07u w=1.6e+07u l=2e+06u
X1 a_2490_n3318# a_2090_n3415# a_2032_n3318# w_n2686_n3537# sky130_fd_pr__pfet_01v8_lvt ad=4.64e+12p pd=3.258e+07u as=4.64e+12p ps=3.258e+07u w=1.6e+07u l=2e+06u
X2 a_n1174_118# a_n1574_21# a_n1632_118# w_n2686_n3537# sky130_fd_pr__pfet_01v8_lvt ad=4.64e+12p pd=3.258e+07u as=0p ps=0u w=1.6e+07u l=2e+06u
X3 a_n258_118# a_n658_21# a_n716_118# w_n2686_n3537# sky130_fd_pr__pfet_01v8_lvt ad=4.64e+12p pd=3.258e+07u as=4.64e+12p ps=3.258e+07u w=1.6e+07u l=2e+06u
X4 a_n716_118# a_n1116_21# a_n1174_118# w_n2686_n3537# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1.6e+07u l=2e+06u
X5 a_1574_n3318# a_1174_n3415# a_1116_n3318# w_n2686_n3537# sky130_fd_pr__pfet_01v8_lvt ad=4.64e+12p pd=3.258e+07u as=4.64e+12p ps=3.258e+07u w=1.6e+07u l=2e+06u
X6 a_n1632_n3318# a_n2032_n3415# a_n2090_n3318# w_n2686_n3537# sky130_fd_pr__pfet_01v8_lvt ad=4.64e+12p pd=3.258e+07u as=4.64e+12p ps=3.258e+07u w=1.6e+07u l=2e+06u
X7 a_n1174_n3318# a_n1574_n3415# a_n1632_n3318# w_n2686_n3537# sky130_fd_pr__pfet_01v8_lvt ad=4.64e+12p pd=3.258e+07u as=0p ps=0u w=1.6e+07u l=2e+06u
X8 a_200_n3318# a_n200_n3415# a_n258_n3318# w_n2686_n3537# sky130_fd_pr__pfet_01v8_lvt ad=4.64e+12p pd=3.258e+07u as=4.64e+12p ps=3.258e+07u w=1.6e+07u l=2e+06u
X9 a_658_118# a_258_21# a_200_118# w_n2686_n3537# sky130_fd_pr__pfet_01v8_lvt ad=4.64e+12p pd=3.258e+07u as=4.64e+12p ps=3.258e+07u w=1.6e+07u l=2e+06u
X10 a_2490_118# a_2090_21# a_2032_118# w_n2686_n3537# sky130_fd_pr__pfet_01v8_lvt ad=4.64e+12p pd=3.258e+07u as=4.64e+12p ps=3.258e+07u w=1.6e+07u l=2e+06u
X11 a_n2090_n3318# a_n2490_n3415# a_n2548_n3318# w_n2686_n3537# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=4.64e+12p ps=3.258e+07u w=1.6e+07u l=2e+06u
X12 a_2032_n3318# a_1632_n3415# a_1574_n3318# w_n2686_n3537# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1.6e+07u l=2e+06u
X13 a_n258_n3318# a_n658_n3415# a_n716_n3318# w_n2686_n3537# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=4.64e+12p ps=3.258e+07u w=1.6e+07u l=2e+06u
X14 a_1116_118# a_716_21# a_658_118# w_n2686_n3537# sky130_fd_pr__pfet_01v8_lvt ad=4.64e+12p pd=3.258e+07u as=0p ps=0u w=1.6e+07u l=2e+06u
X15 a_1574_118# a_1174_21# a_1116_118# w_n2686_n3537# sky130_fd_pr__pfet_01v8_lvt ad=4.64e+12p pd=3.258e+07u as=0p ps=0u w=1.6e+07u l=2e+06u
X16 a_n716_n3318# a_n1116_n3415# a_n1174_n3318# w_n2686_n3537# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1.6e+07u l=2e+06u
X17 a_658_n3318# a_258_n3415# a_200_n3318# w_n2686_n3537# sky130_fd_pr__pfet_01v8_lvt ad=4.64e+12p pd=3.258e+07u as=0p ps=0u w=1.6e+07u l=2e+06u
X18 a_1116_n3318# a_716_n3415# a_658_n3318# w_n2686_n3537# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1.6e+07u l=2e+06u
X19 a_2032_118# a_1632_21# a_1574_118# w_n2686_n3537# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1.6e+07u l=2e+06u
X20 a_200_118# a_n200_21# a_n258_118# w_n2686_n3537# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1.6e+07u l=2e+06u
X21 a_n2090_118# a_n2490_21# a_n2548_118# w_n2686_n3537# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=4.64e+12p ps=3.258e+07u w=1.6e+07u l=2e+06u
.ends

.subckt bias m1_1080_870# m1_1080_160# m1_1510_6800# li_80_4480# VSUBS
Xsky130_fd_pr__nfet_01v8_lvt_J9QE6F_1 VSUBS m1_1080_160# VSUBS m1_1080_160# m1_640_380#
+ VSUBS VSUBS m1_1080_160# VSUBS m1_640_380# VSUBS VSUBS m1_1080_160# m1_640_380#
+ m1_1080_160# m1_640_380# VSUBS m1_1080_160# VSUBS m1_640_380# m1_1080_160# m1_1080_160#
+ VSUBS m1_1080_160# sky130_fd_pr__nfet_01v8_lvt_J9QE6F
Xsky130_fd_pr__pfet_01v8_lvt_QH9SH3_0 li_80_4480# li_80_4480# m1_1070_700# li_80_4480#
+ m1_1070_700# li_80_4480# li_80_4480# m1_1070_700# li_80_4480# m1_1070_700# m1_1070_700#
+ li_80_4480# m1_1510_6800# m1_1070_700# li_80_4480# li_80_4480# li_80_4480# m1_1070_700#
+ li_80_4480# li_80_4480# m1_1070_700# m1_1070_700# m1_1510_6800# m1_1070_700# li_80_4480#
+ li_80_4480# m1_1070_700# m1_1070_700# li_80_4480# m1_1070_700# m1_1070_700# li_80_4480#
+ m1_1070_700# m1_1070_700# m1_1070_700# li_80_4480# li_80_4480# li_80_4480# li_80_4480#
+ li_80_4480# li_80_4480# m1_1510_6800# m1_1070_700# m1_1070_700# m1_1070_700# li_80_4480#
+ m1_1510_6800# sky130_fd_pr__pfet_01v8_lvt_QH9SH3
Xsky130_fd_pr__nfet_01v8_lvt_M93XMJ_0 m1_1080_870# m1_1080_870# VSUBS VSUBS m1_1070_700#
+ m1_1080_870# m1_640_380# VSUBS m1_1070_700# VSUBS m1_1070_700# VSUBS m1_1080_870#
+ m1_1070_700# m1_1080_870# m1_640_380# m1_640_380# m1_1080_870# m1_1070_700# m1_640_380#
+ m1_1080_870# m1_640_380# m1_1080_870# m1_1080_870# sky130_fd_pr__nfet_01v8_lvt_M93XMJ
.ends

.subckt sky130_fd_pr__cap_mim_m3_1_L46JLG m3_n3150_n6250# c1_n3050_n6150#
X0 c1_n3050_n6150# m3_n3150_n6250# sky130_fd_pr__cap_mim_m3_1 l=3e+07u w=3e+07u
X1 c1_n3050_n6150# m3_n3150_n6250# sky130_fd_pr__cap_mim_m3_1 l=3e+07u w=3e+07u
.ends

.subckt rc_model_6cap m1_15830_n15780# VSUBS
Xsky130_fd_pr__nfet_01v8_lvt_Z6RSN3_0 m1_14820_n13900# m1_16920_n14260# VSUBS m1_15830_n15780#
+ sky130_fd_pr__nfet_01v8_lvt_Z6RSN3
Xsky130_fd_pr__nfet_01v8_lvt_Z6RSN3_1 m1_14820_n15340# m1_16920_n14980# VSUBS m1_15830_n15780#
+ sky130_fd_pr__nfet_01v8_lvt_Z6RSN3
Xsky130_fd_pr__nfet_01v8_lvt_Z6RSN3_3 m1_14840_n13120# m1_16920_n13540# VSUBS m1_15830_n15780#
+ sky130_fd_pr__nfet_01v8_lvt_Z6RSN3
Xsky130_fd_pr__nfet_01v8_lvt_Z6RSN3_2 m1_14820_n13900# m1_16920_n13540# VSUBS m1_15830_n15780#
+ sky130_fd_pr__nfet_01v8_lvt_Z6RSN3
Xsky130_fd_pr__nfet_01v8_lvt_Z6RSN3_4 m1_14820_n14620# m1_16920_n14260# VSUBS m1_15830_n15780#
+ sky130_fd_pr__nfet_01v8_lvt_Z6RSN3
Xsky130_fd_pr__nfet_01v8_lvt_Z6RSN3_5 m1_14820_n14620# m1_16920_n14980# VSUBS m1_15830_n15780#
+ sky130_fd_pr__nfet_01v8_lvt_Z6RSN3
Xsky130_fd_pr__nfet_01v8_lvt_Z6RSN3_6 m1_14820_n15340# m1_16920_n15680# VSUBS m1_15830_n15780#
+ sky130_fd_pr__nfet_01v8_lvt_Z6RSN3
Xsky130_fd_pr__nfet_01v8_lvt_Z6RSN3_7 m1_15830_n15780# m1_16920_n15680# VSUBS m1_15830_n15780#
+ sky130_fd_pr__nfet_01v8_lvt_Z6RSN3
Xsky130_fd_pr__res_xhigh_po_5p73_AW8RAB_0 m1_25400_n4800# m1_15000_n11000# VSUBS m1_25400_n12200#
+ m1_25400_400# m1_15000_n3400# m1_15000_1400# VSUBS m1_25400_n12200# m1_25400_n2200#
+ m1_25400_400# m1_15000_n8400# m1_25400_n4800# m1_15000_n6000# m1_15000_n1000# m1_25400_n2200#
+ m1_15000_n8400# m1_14840_n13120# m1_15000_n6000# m1_15000_n1000# m1_15000_1400#
+ m1_25400_n9600# m1_15000_n11000# m1_25400_n7200# m1_25400_n7200# m1_25400_n9600#
+ m1_15000_n3400# sky130_fd_pr__res_xhigh_po_5p73_AW8RAB
Xsky130_fd_pr__cap_mim_m3_1_L46JLG_0 VSUBS m1_15830_n15780# sky130_fd_pr__cap_mim_m3_1_L46JLG
Xsky130_fd_pr__cap_mim_m3_1_LQXKLG_0 VSUBS m1_15830_n15780# sky130_fd_pr__cap_mim_m3_1_LQXKLG
.ends

.subckt and B VDD VSS A Vout
Xsky130_fd_pr__pfet_01v8_TSNZVH_0 m1_280_n300# VDD VDD B sky130_fd_pr__pfet_01v8_TSNZVH
Xsky130_fd_pr__pfet_01v8_TSNZVH_1 m1_280_n300# VDD VDD A sky130_fd_pr__pfet_01v8_TSNZVH
Xinv_0 m1_280_n300# Vout VDD VSS inv
Xsky130_fd_pr__nfet_01v8_Y5UG24_0 VSS B VSS m1_110_n500# sky130_fd_pr__nfet_01v8_Y5UG24
Xsky130_fd_pr__nfet_01v8_Y5UG24_1 m1_110_n500# A VSS m1_280_n300# sky130_fd_pr__nfet_01v8_Y5UG24
.ends

.subckt x2_to_4_decoder D0 D1 D3 D2 A B VDD VSS
Xinv_0 B B_b VDD VSS inv
Xinv_1 A and_3/A VDD VSS inv
Xand_0 B VDD VSS A D3 and
Xand_1 B VDD VSS and_3/A D2 and
Xand_2 B_b VDD VSS A D1 and
Xand_3 B_b VDD VSS and_3/A D0 and
.ends

.subckt cmos_imager_rc_top sh_clk VDD Vb1 Vb0 Vbias Vout A B VSS rst_b_clk
Xrc_model_8cap_0 Vin_3 VSS rc_model_8cap
X3T_0 Vpixel_out rst_b_clk Vin_1 VDD D1 VSS x3T
X3T_1 Vpixel_out rst_b_clk Vin_3 VDD D3 VSS x3T
X3T_2 Vpixel_out rst_b_clk Vin_2 VDD D2 VSS x3T
Xrc_model_4cap_0 Vin_1 VSS rc_model_4cap
Xsample_hold_0 VSS Vcap opamp_realcomp3_usefinger_0/out sh_clk VDD VSS sample_hold
Xcd_output_0 VSS VDD Vout Vcap cd_output
Xopamp_realcomp3_usefinger_0 opamp_realcomp3_usefinger_0/out Vpixel_out Vbias opamp_realcomp3_usefinger_0/out
+ VDD VSS opamp_realcomp3_usefinger
Xcd_current_0 Vb0 Vb1 Vpixel_out VSS cd_current
Xbias_0 Vb1 Vb0 Vout VDD VSS bias
Xrc_model_6cap_0 Vin_2 VSS rc_model_6cap
X2_to_4_decoder_0 2_to_4_decoder_0/D0 D1 D3 D2 A B VDD VSS x2_to_4_decoder
.ends

.subckt sky130_fd_pr__res_xhigh_po_5p73_UZMRKM a_669_10600# a_n3057_n11032# a_n1815_n11032#
+ a_n3057_10600# a_n1815_10600# a_n3187_n11162# a_669_n11032# a_n573_10600# a_n573_n11032#
+ a_1911_n11032# a_1911_10600#
X0 a_n3057_n11032# a_n3057_10600# a_n3187_n11162# sky130_fd_pr__res_xhigh_po_5p73 l=1.06e+08u
X1 a_n573_n11032# a_n573_10600# a_n3187_n11162# sky130_fd_pr__res_xhigh_po_5p73 l=1.06e+08u
X2 a_n1815_n11032# a_n1815_10600# a_n3187_n11162# sky130_fd_pr__res_xhigh_po_5p73 l=1.06e+08u
X3 a_669_n11032# a_669_10600# a_n3187_n11162# sky130_fd_pr__res_xhigh_po_5p73 l=1.06e+08u
X4 a_1911_n11032# a_1911_10600# a_n3187_n11162# sky130_fd_pr__res_xhigh_po_5p73 l=1.06e+08u
.ends

.subckt XM_Rref sky130_fd_pr__res_xhigh_po_5p73_UZMRKM_0/a_1911_n11032# sky130_fd_pr__res_xhigh_po_5p73_UZMRKM_0/a_n3057_10600#
+ VSUBS
Xsky130_fd_pr__res_xhigh_po_5p73_UZMRKM_0 m1_3616_20636# m1_n110_n995# m1_n110_n995#
+ sky130_fd_pr__res_xhigh_po_5p73_UZMRKM_0/a_n3057_10600# m1_1132_20636# VSUBS m1_2374_n995#
+ m1_1132_20636# m1_2374_n995# sky130_fd_pr__res_xhigh_po_5p73_UZMRKM_0/a_1911_n11032#
+ m1_3616_20636# sky130_fd_pr__res_xhigh_po_5p73_UZMRKM
.ends

.subckt sky130_fd_pr__pfet_01v8_lvt_Q24T46 a_n416_n136# a_n616_n162# w_n812_n284#
+ a_358_n136# a_158_n162# a_100_n136# a_n674_n136# a_n158_n136# a_n358_n162# a_616_n136#
+ a_416_n162# a_n100_n162#
X0 a_358_n136# a_158_n162# a_100_n136# w_n812_n284# sky130_fd_pr__pfet_01v8_lvt ad=2.9e+11p pd=2.58e+06u as=2.9e+11p ps=2.58e+06u w=1e+06u l=1e+06u
X1 a_616_n136# a_416_n162# a_358_n136# w_n812_n284# sky130_fd_pr__pfet_01v8_lvt ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=1e+06u
X2 a_100_n136# a_n100_n162# a_n158_n136# w_n812_n284# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=2.9e+11p ps=2.58e+06u w=1e+06u l=1e+06u
X3 a_n416_n136# a_n616_n162# a_n674_n136# w_n812_n284# sky130_fd_pr__pfet_01v8_lvt ad=2.9e+11p pd=2.58e+06u as=2.9e+11p ps=2.58e+06u w=1e+06u l=1e+06u
X4 a_n158_n136# a_n358_n162# a_n416_n136# w_n812_n284# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
.ends

.subckt sky130_fd_pr__pfet_01v8_lvt_MUVY4U a_n616_n161# a_358_n64# a_n674_n64# a_n158_n64#
+ w_n812_n284# a_158_n161# a_n358_n161# a_416_n161# a_n100_n161# a_616_n64# a_100_n64#
+ a_n416_n64#
X0 a_100_n64# a_n100_n161# a_n158_n64# w_n812_n284# sky130_fd_pr__pfet_01v8_lvt ad=2.9e+11p pd=2.58e+06u as=2.9e+11p ps=2.58e+06u w=1e+06u l=1e+06u
X1 a_616_n64# a_416_n161# a_358_n64# w_n812_n284# sky130_fd_pr__pfet_01v8_lvt ad=2.9e+11p pd=2.58e+06u as=2.9e+11p ps=2.58e+06u w=1e+06u l=1e+06u
X2 a_358_n64# a_158_n161# a_100_n64# w_n812_n284# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X3 a_n416_n64# a_n616_n161# a_n674_n64# w_n812_n284# sky130_fd_pr__pfet_01v8_lvt ad=2.9e+11p pd=2.58e+06u as=2.9e+11p ps=2.58e+06u w=1e+06u l=1e+06u
X4 a_n158_n64# a_n358_n161# a_n416_n64# w_n812_n284# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
.ends

.subckt XM_current_gate m1_30_n420# m1_94_n180# li_818_316# m1_30_260#
Xsky130_fd_pr__pfet_01v8_lvt_Q24T46_0 li_818_316# m1_94_n180# li_818_316# m1_30_n420#
+ m1_94_n180# li_818_316# m1_30_n420# m1_30_260# m1_94_n180# li_818_316# m1_94_n180#
+ m1_94_n180# sky130_fd_pr__pfet_01v8_lvt_Q24T46
Xsky130_fd_pr__pfet_01v8_lvt_MUVY4U_0 m1_94_n180# m1_30_260# m1_30_260# m1_30_n420#
+ li_818_316# m1_94_n180# m1_94_n180# m1_94_n180# m1_94_n180# li_818_316# li_818_316#
+ li_818_316# sky130_fd_pr__pfet_01v8_lvt_MUVY4U
.ends

.subckt XM_current_gate_with_dummy XM_current_gate_8/m1_30_260# XM_current_gate_8/m1_30_n420#
+ XM_current_gate_6/m1_30_n420# XM_current_gate_3/m1_94_n180# XM_current_gate_1/m1_94_n180#
+ XM_current_gate_5/m1_30_n420# XM_current_gate_1/m1_30_260# XM_current_gate_3/m1_30_n420#
+ XM_current_gate_6/m1_94_n180# XM_current_gate_7/m1_30_n420# XM_current_gate_2/m1_94_n180#
+ XM_current_gate_2/m1_30_260# XM_current_gate_5/m1_94_n180# XM_current_gate_4/m1_94_n180#
+ XM_current_gate_4/m1_30_260# XM_current_gate_5/m1_30_260# XM_current_gate_0/m1_30_n420#
+ XM_current_gate_7/m1_30_260# XM_current_gate_4/m1_30_n420# XM_current_gate_1/m1_30_n420#
+ XM_current_gate_0/m1_30_260# XM_current_gate_8/m1_94_n180# XM_current_gate_3/m1_30_260#
+ XM_current_gate_0/m1_94_n180# XM_current_gate_6/m1_30_260# XM_current_gate_7/m1_94_n180#
+ XM_current_gate_8/li_818_316# XM_current_gate_2/m1_30_n420#
XXM_current_gate_0 XM_current_gate_0/m1_30_n420# XM_current_gate_0/m1_94_n180# XM_current_gate_8/li_818_316#
+ XM_current_gate_0/m1_30_260# XM_current_gate
XXM_current_gate_1 XM_current_gate_1/m1_30_n420# XM_current_gate_1/m1_94_n180# XM_current_gate_8/li_818_316#
+ XM_current_gate_1/m1_30_260# XM_current_gate
XXM_current_gate_2 XM_current_gate_2/m1_30_n420# XM_current_gate_2/m1_94_n180# XM_current_gate_8/li_818_316#
+ XM_current_gate_2/m1_30_260# XM_current_gate
XXM_current_gate_3 XM_current_gate_3/m1_30_n420# XM_current_gate_3/m1_94_n180# XM_current_gate_8/li_818_316#
+ XM_current_gate_3/m1_30_260# XM_current_gate
XXM_current_gate_4 XM_current_gate_4/m1_30_n420# XM_current_gate_4/m1_94_n180# XM_current_gate_8/li_818_316#
+ XM_current_gate_4/m1_30_260# XM_current_gate
XXM_current_gate_5 XM_current_gate_5/m1_30_n420# XM_current_gate_5/m1_94_n180# XM_current_gate_8/li_818_316#
+ XM_current_gate_5/m1_30_260# XM_current_gate
XXM_current_gate_6 XM_current_gate_6/m1_30_n420# XM_current_gate_6/m1_94_n180# XM_current_gate_8/li_818_316#
+ XM_current_gate_6/m1_30_260# XM_current_gate
XXM_current_gate_7 XM_current_gate_7/m1_30_n420# XM_current_gate_7/m1_94_n180# XM_current_gate_8/li_818_316#
+ XM_current_gate_7/m1_30_260# XM_current_gate
XXM_current_gate_8 XM_current_gate_8/m1_30_n420# XM_current_gate_8/m1_94_n180# XM_current_gate_8/li_818_316#
+ XM_current_gate_8/m1_30_260# XM_current_gate
.ends

.subckt sky130_fd_pr__nfet_01v8_lvt_E2U6GT a_n458_n469# a_n400_n557# a_400_n469# a_n560_n643#
X0 a_400_n469# a_n400_n557# a_n458_n469# a_n560_n643# sky130_fd_pr__nfet_01v8_lvt ad=1.45e+12p pd=1.058e+07u as=1.45e+12p ps=1.058e+07u w=5e+06u l=4e+06u
.ends

.subckt sky130_fd_pr__nfet_01v8_lvt_H8V8HY a_n360_n1143# a_200_n969# a_n200_n1057#
+ a_n258_n969#
X0 a_200_n969# a_n200_n1057# a_n258_n969# a_n360_n1143# sky130_fd_pr__nfet_01v8_lvt ad=2.9e+12p pd=2.058e+07u as=2.9e+12p ps=2.058e+07u w=1e+07u l=2e+06u
.ends

.subckt sky130_fd_pr__res_high_po_1p41_G3LFBQ a_n141_n10832# a_n271_n10962# a_n141_10400#
X0 a_n141_n10832# a_n141_10400# a_n271_n10962# sky130_fd_pr__res_high_po_1p41 l=1.04e+08u
.ends

.subckt sky130_fd_pr__nfet_01v8_lvt_64DJ5N a_n945_n831# a_n487_n831# a_n29_n831# a_887_n831#
+ a_n887_n857# a_429_n831# a_n429_n857# a_487_n857# a_29_n857# VSUBS
X0 a_429_n831# a_29_n857# a_n29_n831# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=2.32e+12p pd=1.658e+07u as=2.32e+12p ps=1.658e+07u w=8e+06u l=2e+06u
X1 a_887_n831# a_487_n857# a_429_n831# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=2.32e+12p pd=1.658e+07u as=0p ps=0u w=8e+06u l=2e+06u
X2 a_n487_n831# a_n887_n857# a_n945_n831# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=2.32e+12p pd=1.658e+07u as=2.32e+12p ps=1.658e+07u w=8e+06u l=2e+06u
X3 a_n29_n831# a_n429_n857# a_n487_n831# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=8e+06u l=2e+06u
.ends

.subckt sky130_fd_pr__nfet_01v8_lvt_64S6GM a_n945_n769# a_n487_n769# a_n887_n857#
+ a_n29_n769# a_887_n769# a_n429_n857# a_487_n857# a_429_n769# a_29_n857# VSUBS
X0 a_429_n769# a_29_n857# a_n29_n769# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=2.32e+12p pd=1.658e+07u as=2.32e+12p ps=1.658e+07u w=8e+06u l=2e+06u
X1 a_887_n769# a_487_n857# a_429_n769# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=2.32e+12p pd=1.658e+07u as=0p ps=0u w=8e+06u l=2e+06u
X2 a_n487_n769# a_n887_n857# a_n945_n769# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=2.32e+12p pd=1.658e+07u as=2.32e+12p ps=1.658e+07u w=8e+06u l=2e+06u
X3 a_n29_n769# a_n429_n857# a_n487_n769# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=8e+06u l=2e+06u
.ends

.subckt XM_output_mirr sky130_fd_pr__nfet_01v8_lvt_64S6GM_1/VSUBS m1_62_n98# m1_62_n3610#
+ m1_n10_n960# m1_n10_n4460# m1_450_n4460#
Xsky130_fd_pr__nfet_01v8_lvt_64DJ5N_0 m1_n10_n960# m1_450_n4460# m1_n10_n960# m1_n10_n960#
+ m1_62_n98# m1_450_n4460# m1_62_n98# m1_62_n98# m1_62_n98# sky130_fd_pr__nfet_01v8_lvt_64S6GM_1/VSUBS
+ sky130_fd_pr__nfet_01v8_lvt_64DJ5N
Xsky130_fd_pr__nfet_01v8_lvt_64DJ5N_1 m1_n10_n4460# m1_450_n4460# m1_n10_n4460# m1_n10_n4460#
+ m1_62_n3610# m1_450_n4460# m1_62_n3610# m1_62_n3610# m1_62_n3610# sky130_fd_pr__nfet_01v8_lvt_64S6GM_1/VSUBS
+ sky130_fd_pr__nfet_01v8_lvt_64DJ5N
Xsky130_fd_pr__nfet_01v8_lvt_64S6GM_0 m1_n10_n960# m1_450_n4460# m1_62_n98# m1_n10_n960#
+ m1_n10_n960# m1_62_n98# m1_62_n98# m1_450_n4460# m1_62_n98# sky130_fd_pr__nfet_01v8_lvt_64S6GM_1/VSUBS
+ sky130_fd_pr__nfet_01v8_lvt_64S6GM
Xsky130_fd_pr__nfet_01v8_lvt_64S6GM_1 m1_n10_n4460# m1_450_n4460# m1_62_n3610# m1_n10_n4460#
+ m1_n10_n4460# m1_62_n3610# m1_62_n3610# m1_450_n4460# m1_62_n3610# sky130_fd_pr__nfet_01v8_lvt_64S6GM_1/VSUBS
+ sky130_fd_pr__nfet_01v8_lvt_64S6GM
.ends

.subckt XM_output_mirr_combined XM_output_mirr_7/m1_450_n4460# XM_output_mirr_7/m1_62_n98#
+ XM_output_mirr_2/m1_n10_n4460# XM_output_mirr_2/m1_62_n98# XM_output_mirr_2/m1_n10_n960#
+ XM_output_mirr_4/m1_n10_n960# XM_output_mirr_7/m1_62_n3610# XM_output_mirr_2/m1_450_n4460#
+ XM_output_mirr_4/m1_62_n98# XM_output_mirr_2/m1_62_n3610# XM_output_mirr_0/m1_450_n4460#
+ XM_output_mirr_5/m1_62_n98# XM_output_mirr_0/m1_62_n98# XM_output_mirr_6/m1_62_n3610#
+ XM_output_mirr_5/m1_n10_n4460# XM_output_mirr_3/m1_n10_n4460# XM_output_mirr_5/m1_62_n3610#
+ XM_output_mirr_6/m1_450_n4460# XM_output_mirr_3/m1_450_n4460# XM_output_mirr_4/m1_450_n4460#
+ XM_output_mirr_7/m1_n10_n960# XM_output_mirr_0/m1_62_n3610# XM_output_mirr_3/m1_62_n98#
+ XM_output_mirr_6/m1_n10_n4460# XM_output_mirr_5/m1_450_n4460# XM_output_mirr_1/m1_450_n4460#
+ XM_output_mirr_1/m1_n10_n960# XM_output_mirr_6/m1_62_n98# XM_output_mirr_3/m1_62_n3610#
+ XM_output_mirr_6/m1_n10_n960# XM_output_mirr_5/m1_n10_n960# XM_output_mirr_7/m1_n10_n4460#
+ XM_output_mirr_1/m1_n10_n4460# XM_output_mirr_1/m1_62_n98# XM_output_mirr_4/m1_62_n3610#
+ XM_output_mirr_4/m1_n10_n4460# XM_output_mirr_0/m1_n10_n960# XM_output_mirr_0/m1_n10_n4460#
+ XM_output_mirr_1/m1_62_n3610# VSUBS XM_output_mirr_3/m1_n10_n960#
XXM_output_mirr_0 VSUBS XM_output_mirr_0/m1_62_n98# XM_output_mirr_0/m1_62_n3610#
+ XM_output_mirr_0/m1_n10_n960# XM_output_mirr_0/m1_n10_n4460# XM_output_mirr_0/m1_450_n4460#
+ XM_output_mirr
XXM_output_mirr_1 VSUBS XM_output_mirr_1/m1_62_n98# XM_output_mirr_1/m1_62_n3610#
+ XM_output_mirr_1/m1_n10_n960# XM_output_mirr_1/m1_n10_n4460# XM_output_mirr_1/m1_450_n4460#
+ XM_output_mirr
XXM_output_mirr_2 VSUBS XM_output_mirr_2/m1_62_n98# XM_output_mirr_2/m1_62_n3610#
+ XM_output_mirr_2/m1_n10_n960# XM_output_mirr_2/m1_n10_n4460# XM_output_mirr_2/m1_450_n4460#
+ XM_output_mirr
XXM_output_mirr_3 VSUBS XM_output_mirr_3/m1_62_n98# XM_output_mirr_3/m1_62_n3610#
+ XM_output_mirr_3/m1_n10_n960# XM_output_mirr_3/m1_n10_n4460# XM_output_mirr_3/m1_450_n4460#
+ XM_output_mirr
XXM_output_mirr_4 VSUBS XM_output_mirr_4/m1_62_n98# XM_output_mirr_4/m1_62_n3610#
+ XM_output_mirr_4/m1_n10_n960# XM_output_mirr_4/m1_n10_n4460# XM_output_mirr_4/m1_450_n4460#
+ XM_output_mirr
XXM_output_mirr_5 VSUBS XM_output_mirr_5/m1_62_n98# XM_output_mirr_5/m1_62_n3610#
+ XM_output_mirr_5/m1_n10_n960# XM_output_mirr_5/m1_n10_n4460# XM_output_mirr_5/m1_450_n4460#
+ XM_output_mirr
XXM_output_mirr_6 VSUBS XM_output_mirr_6/m1_62_n98# XM_output_mirr_6/m1_62_n3610#
+ XM_output_mirr_6/m1_n10_n960# XM_output_mirr_6/m1_n10_n4460# XM_output_mirr_6/m1_450_n4460#
+ XM_output_mirr
XXM_output_mirr_7 VSUBS XM_output_mirr_7/m1_62_n98# XM_output_mirr_7/m1_62_n3610#
+ XM_output_mirr_7/m1_n10_n960# XM_output_mirr_7/m1_n10_n4460# XM_output_mirr_7/m1_450_n4460#
+ XM_output_mirr
.ends

.subckt XM_output_mirr_combined_with_dummy XM_output_mirr_combined_0/XM_output_mirr_5/m1_n10_n960#
+ XM_output_mirr_combined_0/XM_output_mirr_4/m1_n10_n960# XM_output_mirr_combined_0/XM_output_mirr_3/m1_n10_n960#
+ XM_output_mirr_combined_0/XM_output_mirr_7/m1_n10_n960# XM_output_mirr_combined_0/XM_output_mirr_2/m1_n10_n960#
+ m1_300_5420# m1_740_1920# XM_output_mirr_combined_0/XM_output_mirr_6/m1_n10_n960#
+ XM_output_mirr_combined_0/XM_output_mirr_1/m1_n10_n960# m2_300_360# VSUBS
XXM_output_mirr_combined_0 XM_output_mirr_combined_0/XM_output_mirr_7/m1_450_n4460#
+ m1_300_5420# m2_300_360# m1_300_5420# XM_output_mirr_combined_0/XM_output_mirr_2/m1_n10_n960#
+ XM_output_mirr_combined_0/XM_output_mirr_4/m1_n10_n960# m1_740_1920# XM_output_mirr_combined_0/XM_output_mirr_2/m1_450_n4460#
+ m1_300_5420# m1_740_1920# m1_740_1920# m1_300_5420# m1_300_5420# m1_740_1920# m2_300_360#
+ m2_300_360# m1_740_1920# XM_output_mirr_combined_0/XM_output_mirr_6/m1_450_n4460#
+ XM_output_mirr_combined_0/XM_output_mirr_3/m1_450_n4460# XM_output_mirr_combined_0/XM_output_mirr_4/m1_450_n4460#
+ XM_output_mirr_combined_0/XM_output_mirr_7/m1_n10_n960# m1_740_1920# m1_300_5420#
+ m2_300_360# XM_output_mirr_combined_0/XM_output_mirr_5/m1_450_n4460# XM_output_mirr_combined_0/XM_output_mirr_1/m1_450_n4460#
+ XM_output_mirr_combined_0/XM_output_mirr_1/m1_n10_n960# m1_300_5420# m1_740_1920#
+ XM_output_mirr_combined_0/XM_output_mirr_6/m1_n10_n960# XM_output_mirr_combined_0/XM_output_mirr_5/m1_n10_n960#
+ m2_300_360# m2_300_360# m1_300_5420# m1_740_1920# m2_300_360# m1_300_5420# m2_300_360#
+ m1_740_1920# VSUBS XM_output_mirr_combined_0/XM_output_mirr_3/m1_n10_n960# XM_output_mirr_combined
XXM_output_mirr_combined_1 VSUBS VSUBS VSUBS VSUBS VSUBS VSUBS VSUBS VSUBS VSUBS VSUBS
+ VSUBS VSUBS VSUBS VSUBS VSUBS VSUBS VSUBS VSUBS VSUBS VSUBS VSUBS VSUBS VSUBS VSUBS
+ VSUBS VSUBS VSUBS VSUBS VSUBS VSUBS VSUBS VSUBS VSUBS VSUBS VSUBS VSUBS VSUBS VSUBS
+ VSUBS VSUBS VSUBS XM_output_mirr_combined
XXM_output_mirr_combined_2 VSUBS VSUBS VSUBS VSUBS VSUBS VSUBS VSUBS VSUBS VSUBS VSUBS
+ VSUBS VSUBS VSUBS VSUBS VSUBS VSUBS VSUBS VSUBS VSUBS VSUBS VSUBS VSUBS VSUBS VSUBS
+ VSUBS VSUBS VSUBS VSUBS VSUBS VSUBS VSUBS VSUBS VSUBS VSUBS VSUBS VSUBS VSUBS VSUBS
+ VSUBS VSUBS VSUBS XM_output_mirr_combined
XXM_output_mirr_combined_3 VSUBS VSUBS VSUBS VSUBS VSUBS VSUBS VSUBS VSUBS VSUBS VSUBS
+ VSUBS VSUBS VSUBS VSUBS VSUBS VSUBS VSUBS VSUBS VSUBS VSUBS VSUBS VSUBS VSUBS VSUBS
+ VSUBS VSUBS VSUBS VSUBS VSUBS VSUBS VSUBS VSUBS VSUBS VSUBS VSUBS VSUBS VSUBS VSUBS
+ VSUBS VSUBS VSUBS XM_output_mirr_combined
XXM_output_mirr_combined_4 VSUBS VSUBS VSUBS VSUBS VSUBS VSUBS VSUBS VSUBS VSUBS VSUBS
+ VSUBS VSUBS VSUBS VSUBS VSUBS VSUBS VSUBS VSUBS VSUBS VSUBS VSUBS VSUBS VSUBS VSUBS
+ VSUBS VSUBS VSUBS VSUBS VSUBS VSUBS VSUBS VSUBS VSUBS VSUBS VSUBS VSUBS VSUBS VSUBS
+ VSUBS VSUBS VSUBS XM_output_mirr_combined
XXM_output_mirr_combined_5 VSUBS VSUBS VSUBS VSUBS VSUBS VSUBS VSUBS VSUBS VSUBS VSUBS
+ VSUBS VSUBS VSUBS VSUBS VSUBS VSUBS VSUBS VSUBS VSUBS VSUBS VSUBS VSUBS VSUBS VSUBS
+ VSUBS VSUBS VSUBS VSUBS VSUBS VSUBS VSUBS VSUBS VSUBS VSUBS VSUBS VSUBS VSUBS VSUBS
+ VSUBS VSUBS VSUBS XM_output_mirr_combined
XXM_output_mirr_combined_6 VSUBS VSUBS VSUBS VSUBS VSUBS VSUBS VSUBS VSUBS VSUBS VSUBS
+ VSUBS VSUBS VSUBS VSUBS VSUBS VSUBS VSUBS VSUBS VSUBS VSUBS VSUBS VSUBS VSUBS VSUBS
+ VSUBS VSUBS VSUBS VSUBS VSUBS VSUBS VSUBS VSUBS VSUBS VSUBS VSUBS VSUBS VSUBS VSUBS
+ VSUBS VSUBS VSUBS XM_output_mirr_combined
XXM_output_mirr_combined_7 VSUBS VSUBS VSUBS VSUBS VSUBS VSUBS VSUBS VSUBS VSUBS VSUBS
+ VSUBS VSUBS VSUBS VSUBS VSUBS VSUBS VSUBS VSUBS VSUBS VSUBS VSUBS VSUBS VSUBS VSUBS
+ VSUBS VSUBS VSUBS VSUBS VSUBS VSUBS VSUBS VSUBS VSUBS VSUBS VSUBS VSUBS VSUBS VSUBS
+ VSUBS VSUBS VSUBS XM_output_mirr_combined
XXM_output_mirr_combined_8 VSUBS VSUBS VSUBS VSUBS VSUBS VSUBS VSUBS VSUBS VSUBS VSUBS
+ VSUBS VSUBS VSUBS VSUBS VSUBS VSUBS VSUBS VSUBS VSUBS VSUBS VSUBS VSUBS VSUBS VSUBS
+ VSUBS VSUBS VSUBS VSUBS VSUBS VSUBS VSUBS VSUBS VSUBS VSUBS VSUBS VSUBS VSUBS VSUBS
+ VSUBS VSUBS VSUBS XM_output_mirr_combined
.ends

.subckt sky130_fd_pr__res_high_po_1p41_EL7NMZ a_n271_n5562# a_n141_5000# a_n141_n5432#
X0 a_n141_n5432# a_n141_5000# a_n271_n5562# sky130_fd_pr__res_high_po_1p41 l=5e+07u
.ends

.subckt current_ref Iout0 Iout1 Iout2 Iout3 Iout4 Iout5 Iout6 Vbg Vota_bias VDD voutb1
+ voutb2 VSS
XXM_Rref_0 vd4 VSS VSS XM_Rref
XXM_current_gate_with_dummy_0 VDD VDD VDD VDD Vcurrent_gate VDD voutb2 VDD VDD VDD
+ VDD VDD VDD VDD VDD VDD VDD VDD VDD vd4 VDD VDD VDD VDD VDD VDD VDD VDD XM_current_gate_with_dummy
XXM_current_gate_0 Vota_bias Vcurrent_gate VDD Vota_bias_internal XM_current_gate
Xsky130_fd_pr__nfet_01v8_lvt_E2U6GT_0 Vota_bias_internal Vota_bias_internal VSS VSS
+ sky130_fd_pr__nfet_01v8_lvt_E2U6GT
Xsky130_fd_pr__nfet_01v8_lvt_H8V8HY_0 VSS Vota_bias Vota_bias VSS sky130_fd_pr__nfet_01v8_lvt_H8V8HY
Xsky130_fd_pr__res_high_po_1p41_G3LFBQ_0 vd4 VSS m1_27630_n840# sky130_fd_pr__res_high_po_1p41_G3LFBQ
Xopamp_realcomp3_usefinger_0 Vbg vd4 Vota_bias_internal Vcurrent_gate VDD VSS opamp_realcomp3_usefinger
XXM_output_mirr_combined_with_dummy_0 Iout4 Iout3 Iout2 Iout6 Iout1 voutb2 voutb1
+ Iout5 Iout0 VSS VSS XM_output_mirr_combined_with_dummy
Xsky130_fd_pr__res_high_po_1p41_EL7NMZ_0 VSS VSS m1_27630_n840# sky130_fd_pr__res_high_po_1p41_EL7NMZ
.ends

.subckt sky130_fd_pr__diode_pd2nw_05v5_UW3TFX a_n100_n100# w_n238_n238#
D0 a_n100_n100# w_n238_n238# sky130_fd_pr__diode_pd2nw_05v5 pj=4e+06u area=1e+12p
.ends

.subckt diode li_n20_440# m1_100_200#
Xsky130_fd_pr__diode_pd2nw_05v5_UW3TFX_0 m1_100_200# li_n20_440# sky130_fd_pr__diode_pd2nw_05v5_UW3TFX
.ends

.subckt sky130_fd_pr__nfet_01v8_EDB9KC a_n33_n130# a_15_n42# a_n175_n216# a_n73_n42#
X0 a_15_n42# a_n33_n130# a_n73_n42# a_n175_n216# sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=1.218e+11p ps=1.42e+06u w=420000u l=150000u
.ends

.subckt inductor_4 m4_960_n52800# VSUBS
Xsky130_fd_pr__nfet_01v8_EDB9KC_0 VSUBS VSUBS VSUBS VSUBS sky130_fd_pr__nfet_01v8_EDB9KC
.ends

.subckt user_analog_project_wrapper gpio_analog[0] gpio_analog[10] gpio_analog[11]
+ gpio_analog[12] gpio_analog[13] gpio_analog[14] gpio_analog[15] gpio_analog[16]
+ gpio_analog[17] gpio_analog[1] gpio_analog[2] gpio_analog[3] gpio_analog[4] gpio_analog[5]
+ gpio_analog[6] gpio_analog[7] gpio_analog[8] gpio_analog[9] gpio_noesd[0] gpio_noesd[10]
+ gpio_noesd[11] gpio_noesd[12] gpio_noesd[13] gpio_noesd[14] gpio_noesd[15] gpio_noesd[16]
+ gpio_noesd[17] gpio_noesd[1] gpio_noesd[2] gpio_noesd[3] gpio_noesd[4] gpio_noesd[5]
+ gpio_noesd[6] gpio_noesd[7] gpio_noesd[8] gpio_noesd[9] io_analog[0] io_analog[10]
+ io_analog[1] io_analog[2] io_analog[3] io_analog[7] io_analog[8] io_analog[9] io_analog[4]
+ io_analog[5] io_analog[6] io_clamp_high[0] io_clamp_high[1] io_clamp_high[2] io_clamp_low[0]
+ io_clamp_low[1] io_clamp_low[2] io_in[0] io_in[10] io_in[11] io_in[12] io_in[13]
+ io_in[14] io_in[15] io_in[16] io_in[17] io_in[18] io_in[19] io_in[1] io_in[20] io_in[21]
+ io_in[22] io_in[23] io_in[24] io_in[25] io_in[26] io_in[2] io_in[3] io_in[4] io_in[5]
+ io_in[6] io_in[7] io_in[8] io_in[9] io_in_3v3[0] io_in_3v3[10] io_in_3v3[11] io_in_3v3[12]
+ io_in_3v3[13] io_in_3v3[14] io_in_3v3[15] io_in_3v3[16] io_in_3v3[17] io_in_3v3[18]
+ io_in_3v3[19] io_in_3v3[1] io_in_3v3[20] io_in_3v3[21] io_in_3v3[22] io_in_3v3[23]
+ io_in_3v3[24] io_in_3v3[25] io_in_3v3[26] io_in_3v3[2] io_in_3v3[3] io_in_3v3[4]
+ io_in_3v3[5] io_in_3v3[6] io_in_3v3[7] io_in_3v3[8] io_in_3v3[9] io_oeb[0] io_oeb[10]
+ io_oeb[11] io_oeb[12] io_oeb[13] io_oeb[14] io_oeb[15] io_oeb[16] io_oeb[17] io_oeb[18]
+ io_oeb[19] io_oeb[1] io_oeb[20] io_oeb[21] io_oeb[22] io_oeb[23] io_oeb[24] io_oeb[25]
+ io_oeb[26] io_oeb[2] io_oeb[3] io_oeb[4] io_oeb[5] io_oeb[6] io_oeb[7] io_oeb[8]
+ io_oeb[9] io_out[0] io_out[10] io_out[11] io_out[12] io_out[13] io_out[14] io_out[15]
+ io_out[16] io_out[17] io_out[18] io_out[19] io_out[1] io_out[20] io_out[21] io_out[22]
+ io_out[23] io_out[24] io_out[25] io_out[26] io_out[2] io_out[3] io_out[4] io_out[5]
+ io_out[6] io_out[7] io_out[8] io_out[9] la_data_in[0] la_data_in[100] la_data_in[101]
+ la_data_in[102] la_data_in[103] la_data_in[104] la_data_in[105] la_data_in[106]
+ la_data_in[107] la_data_in[108] la_data_in[109] la_data_in[10] la_data_in[110] la_data_in[111]
+ la_data_in[112] la_data_in[113] la_data_in[114] la_data_in[115] la_data_in[116]
+ la_data_in[117] la_data_in[118] la_data_in[119] la_data_in[11] la_data_in[120] la_data_in[121]
+ la_data_in[122] la_data_in[123] la_data_in[124] la_data_in[125] la_data_in[126]
+ la_data_in[127] la_data_in[12] la_data_in[13] la_data_in[14] la_data_in[15] la_data_in[16]
+ la_data_in[17] la_data_in[18] la_data_in[19] la_data_in[1] la_data_in[20] la_data_in[21]
+ la_data_in[22] la_data_in[23] la_data_in[24] la_data_in[25] la_data_in[26] la_data_in[27]
+ la_data_in[28] la_data_in[29] la_data_in[2] la_data_in[30] la_data_in[31] la_data_in[32]
+ la_data_in[33] la_data_in[34] la_data_in[35] la_data_in[36] la_data_in[37] la_data_in[38]
+ la_data_in[39] la_data_in[3] la_data_in[40] la_data_in[41] la_data_in[42] la_data_in[43]
+ la_data_in[44] la_data_in[45] la_data_in[46] la_data_in[47] la_data_in[48] la_data_in[49]
+ la_data_in[4] la_data_in[50] la_data_in[51] la_data_in[52] la_data_in[53] la_data_in[54]
+ la_data_in[55] la_data_in[56] la_data_in[57] la_data_in[58] la_data_in[59] la_data_in[5]
+ la_data_in[60] la_data_in[61] la_data_in[62] la_data_in[63] la_data_in[64] la_data_in[65]
+ la_data_in[66] la_data_in[67] la_data_in[68] la_data_in[69] la_data_in[6] la_data_in[70]
+ la_data_in[71] la_data_in[72] la_data_in[73] la_data_in[74] la_data_in[75] la_data_in[76]
+ la_data_in[77] la_data_in[78] la_data_in[79] la_data_in[7] la_data_in[80] la_data_in[81]
+ la_data_in[82] la_data_in[83] la_data_in[84] la_data_in[85] la_data_in[86] la_data_in[87]
+ la_data_in[88] la_data_in[89] la_data_in[8] la_data_in[90] la_data_in[91] la_data_in[92]
+ la_data_in[93] la_data_in[94] la_data_in[95] la_data_in[96] la_data_in[97] la_data_in[98]
+ la_data_in[99] la_data_in[9] la_data_out[0] la_data_out[100] la_data_out[101] la_data_out[102]
+ la_data_out[103] la_data_out[104] la_data_out[105] la_data_out[106] la_data_out[107]
+ la_data_out[108] la_data_out[109] la_data_out[10] la_data_out[110] la_data_out[111]
+ la_data_out[112] la_data_out[113] la_data_out[114] la_data_out[115] la_data_out[116]
+ la_data_out[117] la_data_out[118] la_data_out[119] la_data_out[11] la_data_out[120]
+ la_data_out[121] la_data_out[122] la_data_out[123] la_data_out[124] la_data_out[125]
+ la_data_out[126] la_data_out[127] la_data_out[12] la_data_out[13] la_data_out[14]
+ la_data_out[15] la_data_out[16] la_data_out[17] la_data_out[18] la_data_out[19]
+ la_data_out[1] la_data_out[20] la_data_out[21] la_data_out[22] la_data_out[23] la_data_out[24]
+ la_data_out[25] la_data_out[26] la_data_out[27] la_data_out[28] la_data_out[29]
+ la_data_out[2] la_data_out[30] la_data_out[31] la_data_out[32] la_data_out[33] la_data_out[34]
+ la_data_out[35] la_data_out[36] la_data_out[37] la_data_out[38] la_data_out[39]
+ la_data_out[3] la_data_out[40] la_data_out[41] la_data_out[42] la_data_out[43] la_data_out[44]
+ la_data_out[45] la_data_out[46] la_data_out[47] la_data_out[48] la_data_out[49]
+ la_data_out[4] la_data_out[50] la_data_out[51] la_data_out[52] la_data_out[53] la_data_out[54]
+ la_data_out[55] la_data_out[56] la_data_out[57] la_data_out[58] la_data_out[59]
+ la_data_out[5] la_data_out[60] la_data_out[61] la_data_out[62] la_data_out[63] la_data_out[64]
+ la_data_out[65] la_data_out[66] la_data_out[67] la_data_out[68] la_data_out[69]
+ la_data_out[6] la_data_out[70] la_data_out[71] la_data_out[72] la_data_out[73] la_data_out[74]
+ la_data_out[75] la_data_out[76] la_data_out[77] la_data_out[78] la_data_out[79]
+ la_data_out[7] la_data_out[80] la_data_out[81] la_data_out[82] la_data_out[83] la_data_out[84]
+ la_data_out[85] la_data_out[86] la_data_out[87] la_data_out[88] la_data_out[89]
+ la_data_out[8] la_data_out[90] la_data_out[91] la_data_out[92] la_data_out[93] la_data_out[94]
+ la_data_out[95] la_data_out[96] la_data_out[97] la_data_out[98] la_data_out[99]
+ la_data_out[9] la_oenb[0] la_oenb[100] la_oenb[101] la_oenb[102] la_oenb[103] la_oenb[104]
+ la_oenb[105] la_oenb[106] la_oenb[107] la_oenb[108] la_oenb[109] la_oenb[10] la_oenb[110]
+ la_oenb[111] la_oenb[112] la_oenb[113] la_oenb[114] la_oenb[115] la_oenb[116] la_oenb[117]
+ la_oenb[118] la_oenb[119] la_oenb[11] la_oenb[120] la_oenb[121] la_oenb[122] la_oenb[123]
+ la_oenb[124] la_oenb[125] la_oenb[126] la_oenb[127] la_oenb[12] la_oenb[13] la_oenb[14]
+ la_oenb[15] la_oenb[16] la_oenb[17] la_oenb[18] la_oenb[19] la_oenb[1] la_oenb[20]
+ la_oenb[21] la_oenb[22] la_oenb[23] la_oenb[24] la_oenb[25] la_oenb[26] la_oenb[27]
+ la_oenb[28] la_oenb[29] la_oenb[2] la_oenb[30] la_oenb[31] la_oenb[32] la_oenb[33]
+ la_oenb[34] la_oenb[35] la_oenb[36] la_oenb[37] la_oenb[38] la_oenb[39] la_oenb[3]
+ la_oenb[40] la_oenb[41] la_oenb[42] la_oenb[43] la_oenb[44] la_oenb[45] la_oenb[46]
+ la_oenb[47] la_oenb[48] la_oenb[49] la_oenb[4] la_oenb[50] la_oenb[51] la_oenb[52]
+ la_oenb[53] la_oenb[54] la_oenb[55] la_oenb[56] la_oenb[57] la_oenb[58] la_oenb[59]
+ la_oenb[5] la_oenb[60] la_oenb[61] la_oenb[62] la_oenb[63] la_oenb[64] la_oenb[65]
+ la_oenb[66] la_oenb[67] la_oenb[68] la_oenb[69] la_oenb[6] la_oenb[70] la_oenb[71]
+ la_oenb[72] la_oenb[73] la_oenb[74] la_oenb[75] la_oenb[76] la_oenb[77] la_oenb[78]
+ la_oenb[79] la_oenb[7] la_oenb[80] la_oenb[81] la_oenb[82] la_oenb[83] la_oenb[84]
+ la_oenb[85] la_oenb[86] la_oenb[87] la_oenb[88] la_oenb[89] la_oenb[8] la_oenb[90]
+ la_oenb[91] la_oenb[92] la_oenb[93] la_oenb[94] la_oenb[95] la_oenb[96] la_oenb[97]
+ la_oenb[98] la_oenb[99] la_oenb[9] user_clock2 user_irq[0] user_irq[1] user_irq[2]
+ vccd1 vccd2 vdda1 vdda2 vssa1 vssa2 vssd1 vssd2 wb_clk_i wb_rst_i wbs_ack_o wbs_adr_i[0]
+ wbs_adr_i[10] wbs_adr_i[11] wbs_adr_i[12] wbs_adr_i[13] wbs_adr_i[14] wbs_adr_i[15]
+ wbs_adr_i[16] wbs_adr_i[17] wbs_adr_i[18] wbs_adr_i[19] wbs_adr_i[1] wbs_adr_i[20]
+ wbs_adr_i[21] wbs_adr_i[22] wbs_adr_i[23] wbs_adr_i[24] wbs_adr_i[25] wbs_adr_i[26]
+ wbs_adr_i[27] wbs_adr_i[28] wbs_adr_i[29] wbs_adr_i[2] wbs_adr_i[30] wbs_adr_i[31]
+ wbs_adr_i[3] wbs_adr_i[4] wbs_adr_i[5] wbs_adr_i[6] wbs_adr_i[7] wbs_adr_i[8] wbs_adr_i[9]
+ wbs_cyc_i wbs_dat_i[0] wbs_dat_i[10] wbs_dat_i[11] wbs_dat_i[12] wbs_dat_i[13] wbs_dat_i[14]
+ wbs_dat_i[15] wbs_dat_i[16] wbs_dat_i[17] wbs_dat_i[18] wbs_dat_i[19] wbs_dat_i[1]
+ wbs_dat_i[20] wbs_dat_i[21] wbs_dat_i[22] wbs_dat_i[23] wbs_dat_i[24] wbs_dat_i[25]
+ wbs_dat_i[26] wbs_dat_i[27] wbs_dat_i[28] wbs_dat_i[29] wbs_dat_i[2] wbs_dat_i[30]
+ wbs_dat_i[31] wbs_dat_i[3] wbs_dat_i[4] wbs_dat_i[5] wbs_dat_i[6] wbs_dat_i[7] wbs_dat_i[8]
+ wbs_dat_i[9] wbs_dat_o[0] wbs_dat_o[10] wbs_dat_o[11] wbs_dat_o[12] wbs_dat_o[13]
+ wbs_dat_o[14] wbs_dat_o[15] wbs_dat_o[16] wbs_dat_o[17] wbs_dat_o[18] wbs_dat_o[19]
+ wbs_dat_o[1] wbs_dat_o[20] wbs_dat_o[21] wbs_dat_o[22] wbs_dat_o[23] wbs_dat_o[24]
+ wbs_dat_o[25] wbs_dat_o[26] wbs_dat_o[27] wbs_dat_o[28] wbs_dat_o[29] wbs_dat_o[2]
+ wbs_dat_o[30] wbs_dat_o[31] wbs_dat_o[3] wbs_dat_o[4] wbs_dat_o[5] wbs_dat_o[6]
+ wbs_dat_o[7] wbs_dat_o[8] wbs_dat_o[9] wbs_sel_i[0] wbs_sel_i[1] wbs_sel_i[2] wbs_sel_i[3]
+ wbs_stb_i wbs_we_i
XVCO-assembly_0 io_in[18] io_in[17] io_in[16] io_in[15] io_in[14] current_ref_0/Iout0
+ vccd2 vccd2 vssa2 VCO-assembly
Xcmos_imager_rc_top_0 io_in[10] vccd2 current_ref_0/voutb2 current_ref_0/voutb1 current_ref_0/Vota_bias
+ io_analog[5] io_in[12] io_in[11] vssa2 io_in[13] cmos_imager_rc_top
Xcurrent_ref_0 current_ref_0/Iout0 io_analog[6] current_ref_0/Iout2 current_ref_0/Iout3
+ current_ref_0/Iout4 current_ref_0/Iout5 current_ref_0/Iout6 io_analog[7] current_ref_0/Vota_bias
+ vccd2 current_ref_0/voutb1 current_ref_0/voutb2 vssa2 current_ref
Xdiode_0 io_analog[1] io_analog[0] diode
Xinductor_4_0 io_in[22] vssa2 inductor_4
.ends

