magic
tech sky130A
magscale 1 2
timestamp 1672327708
<< pwell >>
rect -8191 -5598 8191 5598
<< psubdiff >>
rect -8155 5528 -8059 5562
rect 8059 5528 8155 5562
rect -8155 -5528 -8121 5528
rect 8121 -5528 8155 5528
rect -8155 -5562 -8059 -5528
rect 8059 -5562 8155 -5528
<< psubdiffcont >>
rect -8059 5528 8059 5562
rect -8059 -5562 8059 -5528
<< xpolycontact >>
rect -8025 5000 -6879 5432
rect -8025 -5432 -6879 -5000
rect -6783 5000 -5637 5432
rect -6783 -5432 -5637 -5000
rect -5541 5000 -4395 5432
rect -5541 -5432 -4395 -5000
rect -4299 5000 -3153 5432
rect -4299 -5432 -3153 -5000
rect -3057 5000 -1911 5432
rect -3057 -5432 -1911 -5000
rect -1815 5000 -669 5432
rect -1815 -5432 -669 -5000
rect -573 5000 573 5432
rect -573 -5432 573 -5000
rect 669 5000 1815 5432
rect 669 -5432 1815 -5000
rect 1911 5000 3057 5432
rect 1911 -5432 3057 -5000
rect 3153 5000 4299 5432
rect 3153 -5432 4299 -5000
rect 4395 5000 5541 5432
rect 4395 -5432 5541 -5000
rect 5637 5000 6783 5432
rect 5637 -5432 6783 -5000
rect 6879 5000 8025 5432
rect 6879 -5432 8025 -5000
<< xpolyres >>
rect -8025 -5000 -6879 5000
rect -6783 -5000 -5637 5000
rect -5541 -5000 -4395 5000
rect -4299 -5000 -3153 5000
rect -3057 -5000 -1911 5000
rect -1815 -5000 -669 5000
rect -573 -5000 573 5000
rect 669 -5000 1815 5000
rect 1911 -5000 3057 5000
rect 3153 -5000 4299 5000
rect 4395 -5000 5541 5000
rect 5637 -5000 6783 5000
rect 6879 -5000 8025 5000
<< locali >>
rect -8155 5528 -8059 5562
rect 8059 5528 8155 5562
rect -8155 -5528 -8121 5528
rect 8121 -5528 8155 5528
rect -8155 -5562 -8059 -5528
rect 8059 -5562 8155 -5528
<< viali >>
rect -8009 5017 -6895 5414
rect -6767 5017 -5653 5414
rect -5525 5017 -4411 5414
rect -4283 5017 -3169 5414
rect -3041 5017 -1927 5414
rect -1799 5017 -685 5414
rect -557 5017 557 5414
rect 685 5017 1799 5414
rect 1927 5017 3041 5414
rect 3169 5017 4283 5414
rect 4411 5017 5525 5414
rect 5653 5017 6767 5414
rect 6895 5017 8009 5414
rect -8009 -5414 -6895 -5017
rect -6767 -5414 -5653 -5017
rect -5525 -5414 -4411 -5017
rect -4283 -5414 -3169 -5017
rect -3041 -5414 -1927 -5017
rect -1799 -5414 -685 -5017
rect -557 -5414 557 -5017
rect 685 -5414 1799 -5017
rect 1927 -5414 3041 -5017
rect 3169 -5414 4283 -5017
rect 4411 -5414 5525 -5017
rect 5653 -5414 6767 -5017
rect 6895 -5414 8009 -5017
<< metal1 >>
rect -8021 5414 -6883 5420
rect -8021 5017 -8009 5414
rect -6895 5017 -6883 5414
rect -8021 5011 -6883 5017
rect -6779 5414 -5641 5420
rect -6779 5017 -6767 5414
rect -5653 5017 -5641 5414
rect -6779 5011 -5641 5017
rect -5537 5414 -4399 5420
rect -5537 5017 -5525 5414
rect -4411 5017 -4399 5414
rect -5537 5011 -4399 5017
rect -4295 5414 -3157 5420
rect -4295 5017 -4283 5414
rect -3169 5017 -3157 5414
rect -4295 5011 -3157 5017
rect -3053 5414 -1915 5420
rect -3053 5017 -3041 5414
rect -1927 5017 -1915 5414
rect -3053 5011 -1915 5017
rect -1811 5414 -673 5420
rect -1811 5017 -1799 5414
rect -685 5017 -673 5414
rect -1811 5011 -673 5017
rect -569 5414 569 5420
rect -569 5017 -557 5414
rect 557 5017 569 5414
rect -569 5011 569 5017
rect 673 5414 1811 5420
rect 673 5017 685 5414
rect 1799 5017 1811 5414
rect 673 5011 1811 5017
rect 1915 5414 3053 5420
rect 1915 5017 1927 5414
rect 3041 5017 3053 5414
rect 1915 5011 3053 5017
rect 3157 5414 4295 5420
rect 3157 5017 3169 5414
rect 4283 5017 4295 5414
rect 3157 5011 4295 5017
rect 4399 5414 5537 5420
rect 4399 5017 4411 5414
rect 5525 5017 5537 5414
rect 4399 5011 5537 5017
rect 5641 5414 6779 5420
rect 5641 5017 5653 5414
rect 6767 5017 6779 5414
rect 5641 5011 6779 5017
rect 6883 5414 8021 5420
rect 6883 5017 6895 5414
rect 8009 5017 8021 5414
rect 6883 5011 8021 5017
rect -8021 -5017 -6883 -5011
rect -8021 -5414 -8009 -5017
rect -6895 -5414 -6883 -5017
rect -8021 -5420 -6883 -5414
rect -6779 -5017 -5641 -5011
rect -6779 -5414 -6767 -5017
rect -5653 -5414 -5641 -5017
rect -6779 -5420 -5641 -5414
rect -5537 -5017 -4399 -5011
rect -5537 -5414 -5525 -5017
rect -4411 -5414 -4399 -5017
rect -5537 -5420 -4399 -5414
rect -4295 -5017 -3157 -5011
rect -4295 -5414 -4283 -5017
rect -3169 -5414 -3157 -5017
rect -4295 -5420 -3157 -5414
rect -3053 -5017 -1915 -5011
rect -3053 -5414 -3041 -5017
rect -1927 -5414 -1915 -5017
rect -3053 -5420 -1915 -5414
rect -1811 -5017 -673 -5011
rect -1811 -5414 -1799 -5017
rect -685 -5414 -673 -5017
rect -1811 -5420 -673 -5414
rect -569 -5017 569 -5011
rect -569 -5414 -557 -5017
rect 557 -5414 569 -5017
rect -569 -5420 569 -5414
rect 673 -5017 1811 -5011
rect 673 -5414 685 -5017
rect 1799 -5414 1811 -5017
rect 673 -5420 1811 -5414
rect 1915 -5017 3053 -5011
rect 1915 -5414 1927 -5017
rect 3041 -5414 3053 -5017
rect 1915 -5420 3053 -5414
rect 3157 -5017 4295 -5011
rect 3157 -5414 3169 -5017
rect 4283 -5414 4295 -5017
rect 3157 -5420 4295 -5414
rect 4399 -5017 5537 -5011
rect 4399 -5414 4411 -5017
rect 5525 -5414 5537 -5017
rect 4399 -5420 5537 -5414
rect 5641 -5017 6779 -5011
rect 5641 -5414 5653 -5017
rect 6767 -5414 6779 -5017
rect 5641 -5420 6779 -5414
rect 6883 -5017 8021 -5011
rect 6883 -5414 6895 -5017
rect 8009 -5414 8021 -5017
rect 6883 -5420 8021 -5414
<< res5p73 >>
rect -8027 -5002 -6877 5002
rect -6785 -5002 -5635 5002
rect -5543 -5002 -4393 5002
rect -4301 -5002 -3151 5002
rect -3059 -5002 -1909 5002
rect -1817 -5002 -667 5002
rect -575 -5002 575 5002
rect 667 -5002 1817 5002
rect 1909 -5002 3059 5002
rect 3151 -5002 4301 5002
rect 4393 -5002 5543 5002
rect 5635 -5002 6785 5002
rect 6877 -5002 8027 5002
<< properties >>
string FIXED_BBOX -8138 -5545 8138 5545
string gencell sky130_fd_pr__res_xhigh_po_5p73
string library sky130
string parameters w 5.73 l 50 m 1 nx 13 wmin 5.730 lmin 0.50 rho 2000 val 17.517k dummy 0 dw 0.0 term 188.2 sterm 0.0 caplen 0 wmax 5.730 guard 1 glc 0 grc 0 gtc 1 gbc 1 compatible {sky130_fd_pr__res_xhigh_po_0p35  sky130_fd_pr__res_xhigh_po_0p69 sky130_fd_pr__res_xhigh_po_1p41  sky130_fd_pr__res_xhigh_po_2p85 sky130_fd_pr__res_xhigh_po_5p73} snake 0 full_metal 1 n_guard 0 hv_guard 0 vias 1 viagb 0 viagt 0 viagl 0 viagr 0
<< end >>
