magic
tech sky130A
magscale 1 2
timestamp 1671676230
<< pwell >>
rect -246 -719 246 719
<< nmoslvt >>
rect -50 109 50 509
rect -50 -509 50 -109
<< ndiff >>
rect -108 497 -50 509
rect -108 121 -96 497
rect -62 121 -50 497
rect -108 109 -50 121
rect 50 497 108 509
rect 50 121 62 497
rect 96 121 108 497
rect 50 109 108 121
rect -108 -121 -50 -109
rect -108 -497 -96 -121
rect -62 -497 -50 -121
rect -108 -509 -50 -497
rect 50 -121 108 -109
rect 50 -497 62 -121
rect 96 -497 108 -121
rect 50 -509 108 -497
<< ndiffc >>
rect -96 121 -62 497
rect 62 121 96 497
rect -96 -497 -62 -121
rect 62 -497 96 -121
<< psubdiff >>
rect -210 649 -114 683
rect 114 649 210 683
rect -210 -649 -176 649
rect 176 -649 210 649
rect -210 -683 -114 -649
rect 114 -683 210 -649
<< psubdiffcont >>
rect -114 649 114 683
rect -114 -683 114 -649
<< poly >>
rect -50 581 50 597
rect -50 547 -34 581
rect 34 547 50 581
rect -50 509 50 547
rect -50 71 50 109
rect -50 37 -34 71
rect 34 37 50 71
rect -50 21 50 37
rect -50 -37 50 -21
rect -50 -71 -34 -37
rect 34 -71 50 -37
rect -50 -109 50 -71
rect -50 -547 50 -509
rect -50 -581 -34 -547
rect 34 -581 50 -547
rect -50 -597 50 -581
<< polycont >>
rect -34 547 34 581
rect -34 37 34 71
rect -34 -71 34 -37
rect -34 -581 34 -547
<< locali >>
rect -210 649 -114 683
rect 114 649 210 683
rect -210 -649 -176 649
rect -50 547 -34 581
rect 34 547 50 581
rect -96 497 -62 513
rect -96 105 -62 121
rect 62 497 96 513
rect 62 105 96 121
rect -50 37 -34 71
rect 34 37 50 71
rect -50 -71 -34 -37
rect 34 -71 50 -37
rect -96 -121 -62 -105
rect -96 -513 -62 -497
rect 62 -121 96 -105
rect 62 -513 96 -497
rect -50 -581 -34 -547
rect 34 -581 50 -547
rect 176 -649 210 649
rect -210 -683 -114 -649
rect 114 -683 210 -649
<< viali >>
rect -34 547 34 581
rect -96 121 -62 497
rect 62 121 96 497
rect -34 37 34 71
rect -34 -71 34 -37
rect -96 -497 -62 -121
rect 62 -497 96 -121
rect -34 -581 34 -547
<< metal1 >>
rect -46 581 46 587
rect -46 547 -34 581
rect 34 547 46 581
rect -46 541 46 547
rect -102 497 -56 509
rect -102 121 -96 497
rect -62 121 -56 497
rect -102 109 -56 121
rect 56 497 102 509
rect 56 121 62 497
rect 96 121 102 497
rect 56 109 102 121
rect -46 71 46 77
rect -46 37 -34 71
rect 34 37 46 71
rect -46 31 46 37
rect -46 -37 46 -31
rect -46 -71 -34 -37
rect 34 -71 46 -37
rect -46 -77 46 -71
rect -102 -121 -56 -109
rect -102 -497 -96 -121
rect -62 -497 -56 -121
rect -102 -509 -56 -497
rect 56 -121 102 -109
rect 56 -497 62 -121
rect 96 -497 102 -121
rect 56 -509 102 -497
rect -46 -547 46 -541
rect -46 -581 -34 -547
rect 34 -581 46 -547
rect -46 -587 46 -581
<< properties >>
string FIXED_BBOX -193 -666 193 666
string gencell sky130_fd_pr__nfet_01v8_lvt
string library sky130
string parameters w 2 l 0.5 m 2 nf 1 diffcov 100 polycov 100 guard 1 glc 0 grc 0 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
