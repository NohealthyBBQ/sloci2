magic
tech sky130A
magscale 1 2
timestamp 1662412052
<< error_p >>
rect -8141 172 -8083 178
rect -7949 172 -7891 178
rect -7757 172 -7699 178
rect -7565 172 -7507 178
rect -7373 172 -7315 178
rect -7181 172 -7123 178
rect -6989 172 -6931 178
rect -6797 172 -6739 178
rect -6605 172 -6547 178
rect -6413 172 -6355 178
rect -6221 172 -6163 178
rect -6029 172 -5971 178
rect -5837 172 -5779 178
rect -5645 172 -5587 178
rect -5453 172 -5395 178
rect -5261 172 -5203 178
rect -5069 172 -5011 178
rect -4877 172 -4819 178
rect -4685 172 -4627 178
rect -4493 172 -4435 178
rect -4301 172 -4243 178
rect -4109 172 -4051 178
rect -3917 172 -3859 178
rect -3725 172 -3667 178
rect -3533 172 -3475 178
rect -3341 172 -3283 178
rect -3149 172 -3091 178
rect -2957 172 -2899 178
rect -2765 172 -2707 178
rect -2573 172 -2515 178
rect -2381 172 -2323 178
rect -2189 172 -2131 178
rect -1997 172 -1939 178
rect -1805 172 -1747 178
rect -1613 172 -1555 178
rect -1421 172 -1363 178
rect -1229 172 -1171 178
rect -1037 172 -979 178
rect -845 172 -787 178
rect -653 172 -595 178
rect -461 172 -403 178
rect -269 172 -211 178
rect -77 172 -19 178
rect 115 172 173 178
rect 307 172 365 178
rect 499 172 557 178
rect 691 172 749 178
rect 883 172 941 178
rect 1075 172 1133 178
rect 1267 172 1325 178
rect 1459 172 1517 178
rect 1651 172 1709 178
rect 1843 172 1901 178
rect 2035 172 2093 178
rect 2227 172 2285 178
rect 2419 172 2477 178
rect 2611 172 2669 178
rect 2803 172 2861 178
rect 2995 172 3053 178
rect 3187 172 3245 178
rect 3379 172 3437 178
rect 3571 172 3629 178
rect 3763 172 3821 178
rect 3955 172 4013 178
rect 4147 172 4205 178
rect 4339 172 4397 178
rect 4531 172 4589 178
rect 4723 172 4781 178
rect 4915 172 4973 178
rect 5107 172 5165 178
rect 5299 172 5357 178
rect 5491 172 5549 178
rect 5683 172 5741 178
rect 5875 172 5933 178
rect 6067 172 6125 178
rect 6259 172 6317 178
rect 6451 172 6509 178
rect 6643 172 6701 178
rect 6835 172 6893 178
rect 7027 172 7085 178
rect 7219 172 7277 178
rect 7411 172 7469 178
rect 7603 172 7661 178
rect 7795 172 7853 178
rect 7987 172 8045 178
rect 8179 172 8237 178
rect -8141 138 -8129 172
rect -7949 138 -7937 172
rect -7757 138 -7745 172
rect -7565 138 -7553 172
rect -7373 138 -7361 172
rect -7181 138 -7169 172
rect -6989 138 -6977 172
rect -6797 138 -6785 172
rect -6605 138 -6593 172
rect -6413 138 -6401 172
rect -6221 138 -6209 172
rect -6029 138 -6017 172
rect -5837 138 -5825 172
rect -5645 138 -5633 172
rect -5453 138 -5441 172
rect -5261 138 -5249 172
rect -5069 138 -5057 172
rect -4877 138 -4865 172
rect -4685 138 -4673 172
rect -4493 138 -4481 172
rect -4301 138 -4289 172
rect -4109 138 -4097 172
rect -3917 138 -3905 172
rect -3725 138 -3713 172
rect -3533 138 -3521 172
rect -3341 138 -3329 172
rect -3149 138 -3137 172
rect -2957 138 -2945 172
rect -2765 138 -2753 172
rect -2573 138 -2561 172
rect -2381 138 -2369 172
rect -2189 138 -2177 172
rect -1997 138 -1985 172
rect -1805 138 -1793 172
rect -1613 138 -1601 172
rect -1421 138 -1409 172
rect -1229 138 -1217 172
rect -1037 138 -1025 172
rect -845 138 -833 172
rect -653 138 -641 172
rect -461 138 -449 172
rect -269 138 -257 172
rect -77 138 -65 172
rect 115 138 127 172
rect 307 138 319 172
rect 499 138 511 172
rect 691 138 703 172
rect 883 138 895 172
rect 1075 138 1087 172
rect 1267 138 1279 172
rect 1459 138 1471 172
rect 1651 138 1663 172
rect 1843 138 1855 172
rect 2035 138 2047 172
rect 2227 138 2239 172
rect 2419 138 2431 172
rect 2611 138 2623 172
rect 2803 138 2815 172
rect 2995 138 3007 172
rect 3187 138 3199 172
rect 3379 138 3391 172
rect 3571 138 3583 172
rect 3763 138 3775 172
rect 3955 138 3967 172
rect 4147 138 4159 172
rect 4339 138 4351 172
rect 4531 138 4543 172
rect 4723 138 4735 172
rect 4915 138 4927 172
rect 5107 138 5119 172
rect 5299 138 5311 172
rect 5491 138 5503 172
rect 5683 138 5695 172
rect 5875 138 5887 172
rect 6067 138 6079 172
rect 6259 138 6271 172
rect 6451 138 6463 172
rect 6643 138 6655 172
rect 6835 138 6847 172
rect 7027 138 7039 172
rect 7219 138 7231 172
rect 7411 138 7423 172
rect 7603 138 7615 172
rect 7795 138 7807 172
rect 7987 138 7999 172
rect 8179 138 8191 172
rect -8141 132 -8083 138
rect -7949 132 -7891 138
rect -7757 132 -7699 138
rect -7565 132 -7507 138
rect -7373 132 -7315 138
rect -7181 132 -7123 138
rect -6989 132 -6931 138
rect -6797 132 -6739 138
rect -6605 132 -6547 138
rect -6413 132 -6355 138
rect -6221 132 -6163 138
rect -6029 132 -5971 138
rect -5837 132 -5779 138
rect -5645 132 -5587 138
rect -5453 132 -5395 138
rect -5261 132 -5203 138
rect -5069 132 -5011 138
rect -4877 132 -4819 138
rect -4685 132 -4627 138
rect -4493 132 -4435 138
rect -4301 132 -4243 138
rect -4109 132 -4051 138
rect -3917 132 -3859 138
rect -3725 132 -3667 138
rect -3533 132 -3475 138
rect -3341 132 -3283 138
rect -3149 132 -3091 138
rect -2957 132 -2899 138
rect -2765 132 -2707 138
rect -2573 132 -2515 138
rect -2381 132 -2323 138
rect -2189 132 -2131 138
rect -1997 132 -1939 138
rect -1805 132 -1747 138
rect -1613 132 -1555 138
rect -1421 132 -1363 138
rect -1229 132 -1171 138
rect -1037 132 -979 138
rect -845 132 -787 138
rect -653 132 -595 138
rect -461 132 -403 138
rect -269 132 -211 138
rect -77 132 -19 138
rect 115 132 173 138
rect 307 132 365 138
rect 499 132 557 138
rect 691 132 749 138
rect 883 132 941 138
rect 1075 132 1133 138
rect 1267 132 1325 138
rect 1459 132 1517 138
rect 1651 132 1709 138
rect 1843 132 1901 138
rect 2035 132 2093 138
rect 2227 132 2285 138
rect 2419 132 2477 138
rect 2611 132 2669 138
rect 2803 132 2861 138
rect 2995 132 3053 138
rect 3187 132 3245 138
rect 3379 132 3437 138
rect 3571 132 3629 138
rect 3763 132 3821 138
rect 3955 132 4013 138
rect 4147 132 4205 138
rect 4339 132 4397 138
rect 4531 132 4589 138
rect 4723 132 4781 138
rect 4915 132 4973 138
rect 5107 132 5165 138
rect 5299 132 5357 138
rect 5491 132 5549 138
rect 5683 132 5741 138
rect 5875 132 5933 138
rect 6067 132 6125 138
rect 6259 132 6317 138
rect 6451 132 6509 138
rect 6643 132 6701 138
rect 6835 132 6893 138
rect 7027 132 7085 138
rect 7219 132 7277 138
rect 7411 132 7469 138
rect 7603 132 7661 138
rect 7795 132 7853 138
rect 7987 132 8045 138
rect 8179 132 8237 138
rect -8237 -138 -8179 -132
rect -8045 -138 -7987 -132
rect -7853 -138 -7795 -132
rect -7661 -138 -7603 -132
rect -7469 -138 -7411 -132
rect -7277 -138 -7219 -132
rect -7085 -138 -7027 -132
rect -6893 -138 -6835 -132
rect -6701 -138 -6643 -132
rect -6509 -138 -6451 -132
rect -6317 -138 -6259 -132
rect -6125 -138 -6067 -132
rect -5933 -138 -5875 -132
rect -5741 -138 -5683 -132
rect -5549 -138 -5491 -132
rect -5357 -138 -5299 -132
rect -5165 -138 -5107 -132
rect -4973 -138 -4915 -132
rect -4781 -138 -4723 -132
rect -4589 -138 -4531 -132
rect -4397 -138 -4339 -132
rect -4205 -138 -4147 -132
rect -4013 -138 -3955 -132
rect -3821 -138 -3763 -132
rect -3629 -138 -3571 -132
rect -3437 -138 -3379 -132
rect -3245 -138 -3187 -132
rect -3053 -138 -2995 -132
rect -2861 -138 -2803 -132
rect -2669 -138 -2611 -132
rect -2477 -138 -2419 -132
rect -2285 -138 -2227 -132
rect -2093 -138 -2035 -132
rect -1901 -138 -1843 -132
rect -1709 -138 -1651 -132
rect -1517 -138 -1459 -132
rect -1325 -138 -1267 -132
rect -1133 -138 -1075 -132
rect -941 -138 -883 -132
rect -749 -138 -691 -132
rect -557 -138 -499 -132
rect -365 -138 -307 -132
rect -173 -138 -115 -132
rect 19 -138 77 -132
rect 211 -138 269 -132
rect 403 -138 461 -132
rect 595 -138 653 -132
rect 787 -138 845 -132
rect 979 -138 1037 -132
rect 1171 -138 1229 -132
rect 1363 -138 1421 -132
rect 1555 -138 1613 -132
rect 1747 -138 1805 -132
rect 1939 -138 1997 -132
rect 2131 -138 2189 -132
rect 2323 -138 2381 -132
rect 2515 -138 2573 -132
rect 2707 -138 2765 -132
rect 2899 -138 2957 -132
rect 3091 -138 3149 -132
rect 3283 -138 3341 -132
rect 3475 -138 3533 -132
rect 3667 -138 3725 -132
rect 3859 -138 3917 -132
rect 4051 -138 4109 -132
rect 4243 -138 4301 -132
rect 4435 -138 4493 -132
rect 4627 -138 4685 -132
rect 4819 -138 4877 -132
rect 5011 -138 5069 -132
rect 5203 -138 5261 -132
rect 5395 -138 5453 -132
rect 5587 -138 5645 -132
rect 5779 -138 5837 -132
rect 5971 -138 6029 -132
rect 6163 -138 6221 -132
rect 6355 -138 6413 -132
rect 6547 -138 6605 -132
rect 6739 -138 6797 -132
rect 6931 -138 6989 -132
rect 7123 -138 7181 -132
rect 7315 -138 7373 -132
rect 7507 -138 7565 -132
rect 7699 -138 7757 -132
rect 7891 -138 7949 -132
rect 8083 -138 8141 -132
rect -8237 -172 -8225 -138
rect -8045 -172 -8033 -138
rect -7853 -172 -7841 -138
rect -7661 -172 -7649 -138
rect -7469 -172 -7457 -138
rect -7277 -172 -7265 -138
rect -7085 -172 -7073 -138
rect -6893 -172 -6881 -138
rect -6701 -172 -6689 -138
rect -6509 -172 -6497 -138
rect -6317 -172 -6305 -138
rect -6125 -172 -6113 -138
rect -5933 -172 -5921 -138
rect -5741 -172 -5729 -138
rect -5549 -172 -5537 -138
rect -5357 -172 -5345 -138
rect -5165 -172 -5153 -138
rect -4973 -172 -4961 -138
rect -4781 -172 -4769 -138
rect -4589 -172 -4577 -138
rect -4397 -172 -4385 -138
rect -4205 -172 -4193 -138
rect -4013 -172 -4001 -138
rect -3821 -172 -3809 -138
rect -3629 -172 -3617 -138
rect -3437 -172 -3425 -138
rect -3245 -172 -3233 -138
rect -3053 -172 -3041 -138
rect -2861 -172 -2849 -138
rect -2669 -172 -2657 -138
rect -2477 -172 -2465 -138
rect -2285 -172 -2273 -138
rect -2093 -172 -2081 -138
rect -1901 -172 -1889 -138
rect -1709 -172 -1697 -138
rect -1517 -172 -1505 -138
rect -1325 -172 -1313 -138
rect -1133 -172 -1121 -138
rect -941 -172 -929 -138
rect -749 -172 -737 -138
rect -557 -172 -545 -138
rect -365 -172 -353 -138
rect -173 -172 -161 -138
rect 19 -172 31 -138
rect 211 -172 223 -138
rect 403 -172 415 -138
rect 595 -172 607 -138
rect 787 -172 799 -138
rect 979 -172 991 -138
rect 1171 -172 1183 -138
rect 1363 -172 1375 -138
rect 1555 -172 1567 -138
rect 1747 -172 1759 -138
rect 1939 -172 1951 -138
rect 2131 -172 2143 -138
rect 2323 -172 2335 -138
rect 2515 -172 2527 -138
rect 2707 -172 2719 -138
rect 2899 -172 2911 -138
rect 3091 -172 3103 -138
rect 3283 -172 3295 -138
rect 3475 -172 3487 -138
rect 3667 -172 3679 -138
rect 3859 -172 3871 -138
rect 4051 -172 4063 -138
rect 4243 -172 4255 -138
rect 4435 -172 4447 -138
rect 4627 -172 4639 -138
rect 4819 -172 4831 -138
rect 5011 -172 5023 -138
rect 5203 -172 5215 -138
rect 5395 -172 5407 -138
rect 5587 -172 5599 -138
rect 5779 -172 5791 -138
rect 5971 -172 5983 -138
rect 6163 -172 6175 -138
rect 6355 -172 6367 -138
rect 6547 -172 6559 -138
rect 6739 -172 6751 -138
rect 6931 -172 6943 -138
rect 7123 -172 7135 -138
rect 7315 -172 7327 -138
rect 7507 -172 7519 -138
rect 7699 -172 7711 -138
rect 7891 -172 7903 -138
rect 8083 -172 8095 -138
rect -8237 -178 -8179 -172
rect -8045 -178 -7987 -172
rect -7853 -178 -7795 -172
rect -7661 -178 -7603 -172
rect -7469 -178 -7411 -172
rect -7277 -178 -7219 -172
rect -7085 -178 -7027 -172
rect -6893 -178 -6835 -172
rect -6701 -178 -6643 -172
rect -6509 -178 -6451 -172
rect -6317 -178 -6259 -172
rect -6125 -178 -6067 -172
rect -5933 -178 -5875 -172
rect -5741 -178 -5683 -172
rect -5549 -178 -5491 -172
rect -5357 -178 -5299 -172
rect -5165 -178 -5107 -172
rect -4973 -178 -4915 -172
rect -4781 -178 -4723 -172
rect -4589 -178 -4531 -172
rect -4397 -178 -4339 -172
rect -4205 -178 -4147 -172
rect -4013 -178 -3955 -172
rect -3821 -178 -3763 -172
rect -3629 -178 -3571 -172
rect -3437 -178 -3379 -172
rect -3245 -178 -3187 -172
rect -3053 -178 -2995 -172
rect -2861 -178 -2803 -172
rect -2669 -178 -2611 -172
rect -2477 -178 -2419 -172
rect -2285 -178 -2227 -172
rect -2093 -178 -2035 -172
rect -1901 -178 -1843 -172
rect -1709 -178 -1651 -172
rect -1517 -178 -1459 -172
rect -1325 -178 -1267 -172
rect -1133 -178 -1075 -172
rect -941 -178 -883 -172
rect -749 -178 -691 -172
rect -557 -178 -499 -172
rect -365 -178 -307 -172
rect -173 -178 -115 -172
rect 19 -178 77 -172
rect 211 -178 269 -172
rect 403 -178 461 -172
rect 595 -178 653 -172
rect 787 -178 845 -172
rect 979 -178 1037 -172
rect 1171 -178 1229 -172
rect 1363 -178 1421 -172
rect 1555 -178 1613 -172
rect 1747 -178 1805 -172
rect 1939 -178 1997 -172
rect 2131 -178 2189 -172
rect 2323 -178 2381 -172
rect 2515 -178 2573 -172
rect 2707 -178 2765 -172
rect 2899 -178 2957 -172
rect 3091 -178 3149 -172
rect 3283 -178 3341 -172
rect 3475 -178 3533 -172
rect 3667 -178 3725 -172
rect 3859 -178 3917 -172
rect 4051 -178 4109 -172
rect 4243 -178 4301 -172
rect 4435 -178 4493 -172
rect 4627 -178 4685 -172
rect 4819 -178 4877 -172
rect 5011 -178 5069 -172
rect 5203 -178 5261 -172
rect 5395 -178 5453 -172
rect 5587 -178 5645 -172
rect 5779 -178 5837 -172
rect 5971 -178 6029 -172
rect 6163 -178 6221 -172
rect 6355 -178 6413 -172
rect 6547 -178 6605 -172
rect 6739 -178 6797 -172
rect 6931 -178 6989 -172
rect 7123 -178 7181 -172
rect 7315 -178 7373 -172
rect 7507 -178 7565 -172
rect 7699 -178 7757 -172
rect 7891 -178 7949 -172
rect 8083 -178 8141 -172
<< pwell >>
rect -8423 -310 8423 310
<< nmoslvt >>
rect -8223 -100 -8193 100
rect -8127 -100 -8097 100
rect -8031 -100 -8001 100
rect -7935 -100 -7905 100
rect -7839 -100 -7809 100
rect -7743 -100 -7713 100
rect -7647 -100 -7617 100
rect -7551 -100 -7521 100
rect -7455 -100 -7425 100
rect -7359 -100 -7329 100
rect -7263 -100 -7233 100
rect -7167 -100 -7137 100
rect -7071 -100 -7041 100
rect -6975 -100 -6945 100
rect -6879 -100 -6849 100
rect -6783 -100 -6753 100
rect -6687 -100 -6657 100
rect -6591 -100 -6561 100
rect -6495 -100 -6465 100
rect -6399 -100 -6369 100
rect -6303 -100 -6273 100
rect -6207 -100 -6177 100
rect -6111 -100 -6081 100
rect -6015 -100 -5985 100
rect -5919 -100 -5889 100
rect -5823 -100 -5793 100
rect -5727 -100 -5697 100
rect -5631 -100 -5601 100
rect -5535 -100 -5505 100
rect -5439 -100 -5409 100
rect -5343 -100 -5313 100
rect -5247 -100 -5217 100
rect -5151 -100 -5121 100
rect -5055 -100 -5025 100
rect -4959 -100 -4929 100
rect -4863 -100 -4833 100
rect -4767 -100 -4737 100
rect -4671 -100 -4641 100
rect -4575 -100 -4545 100
rect -4479 -100 -4449 100
rect -4383 -100 -4353 100
rect -4287 -100 -4257 100
rect -4191 -100 -4161 100
rect -4095 -100 -4065 100
rect -3999 -100 -3969 100
rect -3903 -100 -3873 100
rect -3807 -100 -3777 100
rect -3711 -100 -3681 100
rect -3615 -100 -3585 100
rect -3519 -100 -3489 100
rect -3423 -100 -3393 100
rect -3327 -100 -3297 100
rect -3231 -100 -3201 100
rect -3135 -100 -3105 100
rect -3039 -100 -3009 100
rect -2943 -100 -2913 100
rect -2847 -100 -2817 100
rect -2751 -100 -2721 100
rect -2655 -100 -2625 100
rect -2559 -100 -2529 100
rect -2463 -100 -2433 100
rect -2367 -100 -2337 100
rect -2271 -100 -2241 100
rect -2175 -100 -2145 100
rect -2079 -100 -2049 100
rect -1983 -100 -1953 100
rect -1887 -100 -1857 100
rect -1791 -100 -1761 100
rect -1695 -100 -1665 100
rect -1599 -100 -1569 100
rect -1503 -100 -1473 100
rect -1407 -100 -1377 100
rect -1311 -100 -1281 100
rect -1215 -100 -1185 100
rect -1119 -100 -1089 100
rect -1023 -100 -993 100
rect -927 -100 -897 100
rect -831 -100 -801 100
rect -735 -100 -705 100
rect -639 -100 -609 100
rect -543 -100 -513 100
rect -447 -100 -417 100
rect -351 -100 -321 100
rect -255 -100 -225 100
rect -159 -100 -129 100
rect -63 -100 -33 100
rect 33 -100 63 100
rect 129 -100 159 100
rect 225 -100 255 100
rect 321 -100 351 100
rect 417 -100 447 100
rect 513 -100 543 100
rect 609 -100 639 100
rect 705 -100 735 100
rect 801 -100 831 100
rect 897 -100 927 100
rect 993 -100 1023 100
rect 1089 -100 1119 100
rect 1185 -100 1215 100
rect 1281 -100 1311 100
rect 1377 -100 1407 100
rect 1473 -100 1503 100
rect 1569 -100 1599 100
rect 1665 -100 1695 100
rect 1761 -100 1791 100
rect 1857 -100 1887 100
rect 1953 -100 1983 100
rect 2049 -100 2079 100
rect 2145 -100 2175 100
rect 2241 -100 2271 100
rect 2337 -100 2367 100
rect 2433 -100 2463 100
rect 2529 -100 2559 100
rect 2625 -100 2655 100
rect 2721 -100 2751 100
rect 2817 -100 2847 100
rect 2913 -100 2943 100
rect 3009 -100 3039 100
rect 3105 -100 3135 100
rect 3201 -100 3231 100
rect 3297 -100 3327 100
rect 3393 -100 3423 100
rect 3489 -100 3519 100
rect 3585 -100 3615 100
rect 3681 -100 3711 100
rect 3777 -100 3807 100
rect 3873 -100 3903 100
rect 3969 -100 3999 100
rect 4065 -100 4095 100
rect 4161 -100 4191 100
rect 4257 -100 4287 100
rect 4353 -100 4383 100
rect 4449 -100 4479 100
rect 4545 -100 4575 100
rect 4641 -100 4671 100
rect 4737 -100 4767 100
rect 4833 -100 4863 100
rect 4929 -100 4959 100
rect 5025 -100 5055 100
rect 5121 -100 5151 100
rect 5217 -100 5247 100
rect 5313 -100 5343 100
rect 5409 -100 5439 100
rect 5505 -100 5535 100
rect 5601 -100 5631 100
rect 5697 -100 5727 100
rect 5793 -100 5823 100
rect 5889 -100 5919 100
rect 5985 -100 6015 100
rect 6081 -100 6111 100
rect 6177 -100 6207 100
rect 6273 -100 6303 100
rect 6369 -100 6399 100
rect 6465 -100 6495 100
rect 6561 -100 6591 100
rect 6657 -100 6687 100
rect 6753 -100 6783 100
rect 6849 -100 6879 100
rect 6945 -100 6975 100
rect 7041 -100 7071 100
rect 7137 -100 7167 100
rect 7233 -100 7263 100
rect 7329 -100 7359 100
rect 7425 -100 7455 100
rect 7521 -100 7551 100
rect 7617 -100 7647 100
rect 7713 -100 7743 100
rect 7809 -100 7839 100
rect 7905 -100 7935 100
rect 8001 -100 8031 100
rect 8097 -100 8127 100
rect 8193 -100 8223 100
<< ndiff >>
rect -8285 88 -8223 100
rect -8285 -88 -8273 88
rect -8239 -88 -8223 88
rect -8285 -100 -8223 -88
rect -8193 88 -8127 100
rect -8193 -88 -8177 88
rect -8143 -88 -8127 88
rect -8193 -100 -8127 -88
rect -8097 88 -8031 100
rect -8097 -88 -8081 88
rect -8047 -88 -8031 88
rect -8097 -100 -8031 -88
rect -8001 88 -7935 100
rect -8001 -88 -7985 88
rect -7951 -88 -7935 88
rect -8001 -100 -7935 -88
rect -7905 88 -7839 100
rect -7905 -88 -7889 88
rect -7855 -88 -7839 88
rect -7905 -100 -7839 -88
rect -7809 88 -7743 100
rect -7809 -88 -7793 88
rect -7759 -88 -7743 88
rect -7809 -100 -7743 -88
rect -7713 88 -7647 100
rect -7713 -88 -7697 88
rect -7663 -88 -7647 88
rect -7713 -100 -7647 -88
rect -7617 88 -7551 100
rect -7617 -88 -7601 88
rect -7567 -88 -7551 88
rect -7617 -100 -7551 -88
rect -7521 88 -7455 100
rect -7521 -88 -7505 88
rect -7471 -88 -7455 88
rect -7521 -100 -7455 -88
rect -7425 88 -7359 100
rect -7425 -88 -7409 88
rect -7375 -88 -7359 88
rect -7425 -100 -7359 -88
rect -7329 88 -7263 100
rect -7329 -88 -7313 88
rect -7279 -88 -7263 88
rect -7329 -100 -7263 -88
rect -7233 88 -7167 100
rect -7233 -88 -7217 88
rect -7183 -88 -7167 88
rect -7233 -100 -7167 -88
rect -7137 88 -7071 100
rect -7137 -88 -7121 88
rect -7087 -88 -7071 88
rect -7137 -100 -7071 -88
rect -7041 88 -6975 100
rect -7041 -88 -7025 88
rect -6991 -88 -6975 88
rect -7041 -100 -6975 -88
rect -6945 88 -6879 100
rect -6945 -88 -6929 88
rect -6895 -88 -6879 88
rect -6945 -100 -6879 -88
rect -6849 88 -6783 100
rect -6849 -88 -6833 88
rect -6799 -88 -6783 88
rect -6849 -100 -6783 -88
rect -6753 88 -6687 100
rect -6753 -88 -6737 88
rect -6703 -88 -6687 88
rect -6753 -100 -6687 -88
rect -6657 88 -6591 100
rect -6657 -88 -6641 88
rect -6607 -88 -6591 88
rect -6657 -100 -6591 -88
rect -6561 88 -6495 100
rect -6561 -88 -6545 88
rect -6511 -88 -6495 88
rect -6561 -100 -6495 -88
rect -6465 88 -6399 100
rect -6465 -88 -6449 88
rect -6415 -88 -6399 88
rect -6465 -100 -6399 -88
rect -6369 88 -6303 100
rect -6369 -88 -6353 88
rect -6319 -88 -6303 88
rect -6369 -100 -6303 -88
rect -6273 88 -6207 100
rect -6273 -88 -6257 88
rect -6223 -88 -6207 88
rect -6273 -100 -6207 -88
rect -6177 88 -6111 100
rect -6177 -88 -6161 88
rect -6127 -88 -6111 88
rect -6177 -100 -6111 -88
rect -6081 88 -6015 100
rect -6081 -88 -6065 88
rect -6031 -88 -6015 88
rect -6081 -100 -6015 -88
rect -5985 88 -5919 100
rect -5985 -88 -5969 88
rect -5935 -88 -5919 88
rect -5985 -100 -5919 -88
rect -5889 88 -5823 100
rect -5889 -88 -5873 88
rect -5839 -88 -5823 88
rect -5889 -100 -5823 -88
rect -5793 88 -5727 100
rect -5793 -88 -5777 88
rect -5743 -88 -5727 88
rect -5793 -100 -5727 -88
rect -5697 88 -5631 100
rect -5697 -88 -5681 88
rect -5647 -88 -5631 88
rect -5697 -100 -5631 -88
rect -5601 88 -5535 100
rect -5601 -88 -5585 88
rect -5551 -88 -5535 88
rect -5601 -100 -5535 -88
rect -5505 88 -5439 100
rect -5505 -88 -5489 88
rect -5455 -88 -5439 88
rect -5505 -100 -5439 -88
rect -5409 88 -5343 100
rect -5409 -88 -5393 88
rect -5359 -88 -5343 88
rect -5409 -100 -5343 -88
rect -5313 88 -5247 100
rect -5313 -88 -5297 88
rect -5263 -88 -5247 88
rect -5313 -100 -5247 -88
rect -5217 88 -5151 100
rect -5217 -88 -5201 88
rect -5167 -88 -5151 88
rect -5217 -100 -5151 -88
rect -5121 88 -5055 100
rect -5121 -88 -5105 88
rect -5071 -88 -5055 88
rect -5121 -100 -5055 -88
rect -5025 88 -4959 100
rect -5025 -88 -5009 88
rect -4975 -88 -4959 88
rect -5025 -100 -4959 -88
rect -4929 88 -4863 100
rect -4929 -88 -4913 88
rect -4879 -88 -4863 88
rect -4929 -100 -4863 -88
rect -4833 88 -4767 100
rect -4833 -88 -4817 88
rect -4783 -88 -4767 88
rect -4833 -100 -4767 -88
rect -4737 88 -4671 100
rect -4737 -88 -4721 88
rect -4687 -88 -4671 88
rect -4737 -100 -4671 -88
rect -4641 88 -4575 100
rect -4641 -88 -4625 88
rect -4591 -88 -4575 88
rect -4641 -100 -4575 -88
rect -4545 88 -4479 100
rect -4545 -88 -4529 88
rect -4495 -88 -4479 88
rect -4545 -100 -4479 -88
rect -4449 88 -4383 100
rect -4449 -88 -4433 88
rect -4399 -88 -4383 88
rect -4449 -100 -4383 -88
rect -4353 88 -4287 100
rect -4353 -88 -4337 88
rect -4303 -88 -4287 88
rect -4353 -100 -4287 -88
rect -4257 88 -4191 100
rect -4257 -88 -4241 88
rect -4207 -88 -4191 88
rect -4257 -100 -4191 -88
rect -4161 88 -4095 100
rect -4161 -88 -4145 88
rect -4111 -88 -4095 88
rect -4161 -100 -4095 -88
rect -4065 88 -3999 100
rect -4065 -88 -4049 88
rect -4015 -88 -3999 88
rect -4065 -100 -3999 -88
rect -3969 88 -3903 100
rect -3969 -88 -3953 88
rect -3919 -88 -3903 88
rect -3969 -100 -3903 -88
rect -3873 88 -3807 100
rect -3873 -88 -3857 88
rect -3823 -88 -3807 88
rect -3873 -100 -3807 -88
rect -3777 88 -3711 100
rect -3777 -88 -3761 88
rect -3727 -88 -3711 88
rect -3777 -100 -3711 -88
rect -3681 88 -3615 100
rect -3681 -88 -3665 88
rect -3631 -88 -3615 88
rect -3681 -100 -3615 -88
rect -3585 88 -3519 100
rect -3585 -88 -3569 88
rect -3535 -88 -3519 88
rect -3585 -100 -3519 -88
rect -3489 88 -3423 100
rect -3489 -88 -3473 88
rect -3439 -88 -3423 88
rect -3489 -100 -3423 -88
rect -3393 88 -3327 100
rect -3393 -88 -3377 88
rect -3343 -88 -3327 88
rect -3393 -100 -3327 -88
rect -3297 88 -3231 100
rect -3297 -88 -3281 88
rect -3247 -88 -3231 88
rect -3297 -100 -3231 -88
rect -3201 88 -3135 100
rect -3201 -88 -3185 88
rect -3151 -88 -3135 88
rect -3201 -100 -3135 -88
rect -3105 88 -3039 100
rect -3105 -88 -3089 88
rect -3055 -88 -3039 88
rect -3105 -100 -3039 -88
rect -3009 88 -2943 100
rect -3009 -88 -2993 88
rect -2959 -88 -2943 88
rect -3009 -100 -2943 -88
rect -2913 88 -2847 100
rect -2913 -88 -2897 88
rect -2863 -88 -2847 88
rect -2913 -100 -2847 -88
rect -2817 88 -2751 100
rect -2817 -88 -2801 88
rect -2767 -88 -2751 88
rect -2817 -100 -2751 -88
rect -2721 88 -2655 100
rect -2721 -88 -2705 88
rect -2671 -88 -2655 88
rect -2721 -100 -2655 -88
rect -2625 88 -2559 100
rect -2625 -88 -2609 88
rect -2575 -88 -2559 88
rect -2625 -100 -2559 -88
rect -2529 88 -2463 100
rect -2529 -88 -2513 88
rect -2479 -88 -2463 88
rect -2529 -100 -2463 -88
rect -2433 88 -2367 100
rect -2433 -88 -2417 88
rect -2383 -88 -2367 88
rect -2433 -100 -2367 -88
rect -2337 88 -2271 100
rect -2337 -88 -2321 88
rect -2287 -88 -2271 88
rect -2337 -100 -2271 -88
rect -2241 88 -2175 100
rect -2241 -88 -2225 88
rect -2191 -88 -2175 88
rect -2241 -100 -2175 -88
rect -2145 88 -2079 100
rect -2145 -88 -2129 88
rect -2095 -88 -2079 88
rect -2145 -100 -2079 -88
rect -2049 88 -1983 100
rect -2049 -88 -2033 88
rect -1999 -88 -1983 88
rect -2049 -100 -1983 -88
rect -1953 88 -1887 100
rect -1953 -88 -1937 88
rect -1903 -88 -1887 88
rect -1953 -100 -1887 -88
rect -1857 88 -1791 100
rect -1857 -88 -1841 88
rect -1807 -88 -1791 88
rect -1857 -100 -1791 -88
rect -1761 88 -1695 100
rect -1761 -88 -1745 88
rect -1711 -88 -1695 88
rect -1761 -100 -1695 -88
rect -1665 88 -1599 100
rect -1665 -88 -1649 88
rect -1615 -88 -1599 88
rect -1665 -100 -1599 -88
rect -1569 88 -1503 100
rect -1569 -88 -1553 88
rect -1519 -88 -1503 88
rect -1569 -100 -1503 -88
rect -1473 88 -1407 100
rect -1473 -88 -1457 88
rect -1423 -88 -1407 88
rect -1473 -100 -1407 -88
rect -1377 88 -1311 100
rect -1377 -88 -1361 88
rect -1327 -88 -1311 88
rect -1377 -100 -1311 -88
rect -1281 88 -1215 100
rect -1281 -88 -1265 88
rect -1231 -88 -1215 88
rect -1281 -100 -1215 -88
rect -1185 88 -1119 100
rect -1185 -88 -1169 88
rect -1135 -88 -1119 88
rect -1185 -100 -1119 -88
rect -1089 88 -1023 100
rect -1089 -88 -1073 88
rect -1039 -88 -1023 88
rect -1089 -100 -1023 -88
rect -993 88 -927 100
rect -993 -88 -977 88
rect -943 -88 -927 88
rect -993 -100 -927 -88
rect -897 88 -831 100
rect -897 -88 -881 88
rect -847 -88 -831 88
rect -897 -100 -831 -88
rect -801 88 -735 100
rect -801 -88 -785 88
rect -751 -88 -735 88
rect -801 -100 -735 -88
rect -705 88 -639 100
rect -705 -88 -689 88
rect -655 -88 -639 88
rect -705 -100 -639 -88
rect -609 88 -543 100
rect -609 -88 -593 88
rect -559 -88 -543 88
rect -609 -100 -543 -88
rect -513 88 -447 100
rect -513 -88 -497 88
rect -463 -88 -447 88
rect -513 -100 -447 -88
rect -417 88 -351 100
rect -417 -88 -401 88
rect -367 -88 -351 88
rect -417 -100 -351 -88
rect -321 88 -255 100
rect -321 -88 -305 88
rect -271 -88 -255 88
rect -321 -100 -255 -88
rect -225 88 -159 100
rect -225 -88 -209 88
rect -175 -88 -159 88
rect -225 -100 -159 -88
rect -129 88 -63 100
rect -129 -88 -113 88
rect -79 -88 -63 88
rect -129 -100 -63 -88
rect -33 88 33 100
rect -33 -88 -17 88
rect 17 -88 33 88
rect -33 -100 33 -88
rect 63 88 129 100
rect 63 -88 79 88
rect 113 -88 129 88
rect 63 -100 129 -88
rect 159 88 225 100
rect 159 -88 175 88
rect 209 -88 225 88
rect 159 -100 225 -88
rect 255 88 321 100
rect 255 -88 271 88
rect 305 -88 321 88
rect 255 -100 321 -88
rect 351 88 417 100
rect 351 -88 367 88
rect 401 -88 417 88
rect 351 -100 417 -88
rect 447 88 513 100
rect 447 -88 463 88
rect 497 -88 513 88
rect 447 -100 513 -88
rect 543 88 609 100
rect 543 -88 559 88
rect 593 -88 609 88
rect 543 -100 609 -88
rect 639 88 705 100
rect 639 -88 655 88
rect 689 -88 705 88
rect 639 -100 705 -88
rect 735 88 801 100
rect 735 -88 751 88
rect 785 -88 801 88
rect 735 -100 801 -88
rect 831 88 897 100
rect 831 -88 847 88
rect 881 -88 897 88
rect 831 -100 897 -88
rect 927 88 993 100
rect 927 -88 943 88
rect 977 -88 993 88
rect 927 -100 993 -88
rect 1023 88 1089 100
rect 1023 -88 1039 88
rect 1073 -88 1089 88
rect 1023 -100 1089 -88
rect 1119 88 1185 100
rect 1119 -88 1135 88
rect 1169 -88 1185 88
rect 1119 -100 1185 -88
rect 1215 88 1281 100
rect 1215 -88 1231 88
rect 1265 -88 1281 88
rect 1215 -100 1281 -88
rect 1311 88 1377 100
rect 1311 -88 1327 88
rect 1361 -88 1377 88
rect 1311 -100 1377 -88
rect 1407 88 1473 100
rect 1407 -88 1423 88
rect 1457 -88 1473 88
rect 1407 -100 1473 -88
rect 1503 88 1569 100
rect 1503 -88 1519 88
rect 1553 -88 1569 88
rect 1503 -100 1569 -88
rect 1599 88 1665 100
rect 1599 -88 1615 88
rect 1649 -88 1665 88
rect 1599 -100 1665 -88
rect 1695 88 1761 100
rect 1695 -88 1711 88
rect 1745 -88 1761 88
rect 1695 -100 1761 -88
rect 1791 88 1857 100
rect 1791 -88 1807 88
rect 1841 -88 1857 88
rect 1791 -100 1857 -88
rect 1887 88 1953 100
rect 1887 -88 1903 88
rect 1937 -88 1953 88
rect 1887 -100 1953 -88
rect 1983 88 2049 100
rect 1983 -88 1999 88
rect 2033 -88 2049 88
rect 1983 -100 2049 -88
rect 2079 88 2145 100
rect 2079 -88 2095 88
rect 2129 -88 2145 88
rect 2079 -100 2145 -88
rect 2175 88 2241 100
rect 2175 -88 2191 88
rect 2225 -88 2241 88
rect 2175 -100 2241 -88
rect 2271 88 2337 100
rect 2271 -88 2287 88
rect 2321 -88 2337 88
rect 2271 -100 2337 -88
rect 2367 88 2433 100
rect 2367 -88 2383 88
rect 2417 -88 2433 88
rect 2367 -100 2433 -88
rect 2463 88 2529 100
rect 2463 -88 2479 88
rect 2513 -88 2529 88
rect 2463 -100 2529 -88
rect 2559 88 2625 100
rect 2559 -88 2575 88
rect 2609 -88 2625 88
rect 2559 -100 2625 -88
rect 2655 88 2721 100
rect 2655 -88 2671 88
rect 2705 -88 2721 88
rect 2655 -100 2721 -88
rect 2751 88 2817 100
rect 2751 -88 2767 88
rect 2801 -88 2817 88
rect 2751 -100 2817 -88
rect 2847 88 2913 100
rect 2847 -88 2863 88
rect 2897 -88 2913 88
rect 2847 -100 2913 -88
rect 2943 88 3009 100
rect 2943 -88 2959 88
rect 2993 -88 3009 88
rect 2943 -100 3009 -88
rect 3039 88 3105 100
rect 3039 -88 3055 88
rect 3089 -88 3105 88
rect 3039 -100 3105 -88
rect 3135 88 3201 100
rect 3135 -88 3151 88
rect 3185 -88 3201 88
rect 3135 -100 3201 -88
rect 3231 88 3297 100
rect 3231 -88 3247 88
rect 3281 -88 3297 88
rect 3231 -100 3297 -88
rect 3327 88 3393 100
rect 3327 -88 3343 88
rect 3377 -88 3393 88
rect 3327 -100 3393 -88
rect 3423 88 3489 100
rect 3423 -88 3439 88
rect 3473 -88 3489 88
rect 3423 -100 3489 -88
rect 3519 88 3585 100
rect 3519 -88 3535 88
rect 3569 -88 3585 88
rect 3519 -100 3585 -88
rect 3615 88 3681 100
rect 3615 -88 3631 88
rect 3665 -88 3681 88
rect 3615 -100 3681 -88
rect 3711 88 3777 100
rect 3711 -88 3727 88
rect 3761 -88 3777 88
rect 3711 -100 3777 -88
rect 3807 88 3873 100
rect 3807 -88 3823 88
rect 3857 -88 3873 88
rect 3807 -100 3873 -88
rect 3903 88 3969 100
rect 3903 -88 3919 88
rect 3953 -88 3969 88
rect 3903 -100 3969 -88
rect 3999 88 4065 100
rect 3999 -88 4015 88
rect 4049 -88 4065 88
rect 3999 -100 4065 -88
rect 4095 88 4161 100
rect 4095 -88 4111 88
rect 4145 -88 4161 88
rect 4095 -100 4161 -88
rect 4191 88 4257 100
rect 4191 -88 4207 88
rect 4241 -88 4257 88
rect 4191 -100 4257 -88
rect 4287 88 4353 100
rect 4287 -88 4303 88
rect 4337 -88 4353 88
rect 4287 -100 4353 -88
rect 4383 88 4449 100
rect 4383 -88 4399 88
rect 4433 -88 4449 88
rect 4383 -100 4449 -88
rect 4479 88 4545 100
rect 4479 -88 4495 88
rect 4529 -88 4545 88
rect 4479 -100 4545 -88
rect 4575 88 4641 100
rect 4575 -88 4591 88
rect 4625 -88 4641 88
rect 4575 -100 4641 -88
rect 4671 88 4737 100
rect 4671 -88 4687 88
rect 4721 -88 4737 88
rect 4671 -100 4737 -88
rect 4767 88 4833 100
rect 4767 -88 4783 88
rect 4817 -88 4833 88
rect 4767 -100 4833 -88
rect 4863 88 4929 100
rect 4863 -88 4879 88
rect 4913 -88 4929 88
rect 4863 -100 4929 -88
rect 4959 88 5025 100
rect 4959 -88 4975 88
rect 5009 -88 5025 88
rect 4959 -100 5025 -88
rect 5055 88 5121 100
rect 5055 -88 5071 88
rect 5105 -88 5121 88
rect 5055 -100 5121 -88
rect 5151 88 5217 100
rect 5151 -88 5167 88
rect 5201 -88 5217 88
rect 5151 -100 5217 -88
rect 5247 88 5313 100
rect 5247 -88 5263 88
rect 5297 -88 5313 88
rect 5247 -100 5313 -88
rect 5343 88 5409 100
rect 5343 -88 5359 88
rect 5393 -88 5409 88
rect 5343 -100 5409 -88
rect 5439 88 5505 100
rect 5439 -88 5455 88
rect 5489 -88 5505 88
rect 5439 -100 5505 -88
rect 5535 88 5601 100
rect 5535 -88 5551 88
rect 5585 -88 5601 88
rect 5535 -100 5601 -88
rect 5631 88 5697 100
rect 5631 -88 5647 88
rect 5681 -88 5697 88
rect 5631 -100 5697 -88
rect 5727 88 5793 100
rect 5727 -88 5743 88
rect 5777 -88 5793 88
rect 5727 -100 5793 -88
rect 5823 88 5889 100
rect 5823 -88 5839 88
rect 5873 -88 5889 88
rect 5823 -100 5889 -88
rect 5919 88 5985 100
rect 5919 -88 5935 88
rect 5969 -88 5985 88
rect 5919 -100 5985 -88
rect 6015 88 6081 100
rect 6015 -88 6031 88
rect 6065 -88 6081 88
rect 6015 -100 6081 -88
rect 6111 88 6177 100
rect 6111 -88 6127 88
rect 6161 -88 6177 88
rect 6111 -100 6177 -88
rect 6207 88 6273 100
rect 6207 -88 6223 88
rect 6257 -88 6273 88
rect 6207 -100 6273 -88
rect 6303 88 6369 100
rect 6303 -88 6319 88
rect 6353 -88 6369 88
rect 6303 -100 6369 -88
rect 6399 88 6465 100
rect 6399 -88 6415 88
rect 6449 -88 6465 88
rect 6399 -100 6465 -88
rect 6495 88 6561 100
rect 6495 -88 6511 88
rect 6545 -88 6561 88
rect 6495 -100 6561 -88
rect 6591 88 6657 100
rect 6591 -88 6607 88
rect 6641 -88 6657 88
rect 6591 -100 6657 -88
rect 6687 88 6753 100
rect 6687 -88 6703 88
rect 6737 -88 6753 88
rect 6687 -100 6753 -88
rect 6783 88 6849 100
rect 6783 -88 6799 88
rect 6833 -88 6849 88
rect 6783 -100 6849 -88
rect 6879 88 6945 100
rect 6879 -88 6895 88
rect 6929 -88 6945 88
rect 6879 -100 6945 -88
rect 6975 88 7041 100
rect 6975 -88 6991 88
rect 7025 -88 7041 88
rect 6975 -100 7041 -88
rect 7071 88 7137 100
rect 7071 -88 7087 88
rect 7121 -88 7137 88
rect 7071 -100 7137 -88
rect 7167 88 7233 100
rect 7167 -88 7183 88
rect 7217 -88 7233 88
rect 7167 -100 7233 -88
rect 7263 88 7329 100
rect 7263 -88 7279 88
rect 7313 -88 7329 88
rect 7263 -100 7329 -88
rect 7359 88 7425 100
rect 7359 -88 7375 88
rect 7409 -88 7425 88
rect 7359 -100 7425 -88
rect 7455 88 7521 100
rect 7455 -88 7471 88
rect 7505 -88 7521 88
rect 7455 -100 7521 -88
rect 7551 88 7617 100
rect 7551 -88 7567 88
rect 7601 -88 7617 88
rect 7551 -100 7617 -88
rect 7647 88 7713 100
rect 7647 -88 7663 88
rect 7697 -88 7713 88
rect 7647 -100 7713 -88
rect 7743 88 7809 100
rect 7743 -88 7759 88
rect 7793 -88 7809 88
rect 7743 -100 7809 -88
rect 7839 88 7905 100
rect 7839 -88 7855 88
rect 7889 -88 7905 88
rect 7839 -100 7905 -88
rect 7935 88 8001 100
rect 7935 -88 7951 88
rect 7985 -88 8001 88
rect 7935 -100 8001 -88
rect 8031 88 8097 100
rect 8031 -88 8047 88
rect 8081 -88 8097 88
rect 8031 -100 8097 -88
rect 8127 88 8193 100
rect 8127 -88 8143 88
rect 8177 -88 8193 88
rect 8127 -100 8193 -88
rect 8223 88 8285 100
rect 8223 -88 8239 88
rect 8273 -88 8285 88
rect 8223 -100 8285 -88
<< ndiffc >>
rect -8273 -88 -8239 88
rect -8177 -88 -8143 88
rect -8081 -88 -8047 88
rect -7985 -88 -7951 88
rect -7889 -88 -7855 88
rect -7793 -88 -7759 88
rect -7697 -88 -7663 88
rect -7601 -88 -7567 88
rect -7505 -88 -7471 88
rect -7409 -88 -7375 88
rect -7313 -88 -7279 88
rect -7217 -88 -7183 88
rect -7121 -88 -7087 88
rect -7025 -88 -6991 88
rect -6929 -88 -6895 88
rect -6833 -88 -6799 88
rect -6737 -88 -6703 88
rect -6641 -88 -6607 88
rect -6545 -88 -6511 88
rect -6449 -88 -6415 88
rect -6353 -88 -6319 88
rect -6257 -88 -6223 88
rect -6161 -88 -6127 88
rect -6065 -88 -6031 88
rect -5969 -88 -5935 88
rect -5873 -88 -5839 88
rect -5777 -88 -5743 88
rect -5681 -88 -5647 88
rect -5585 -88 -5551 88
rect -5489 -88 -5455 88
rect -5393 -88 -5359 88
rect -5297 -88 -5263 88
rect -5201 -88 -5167 88
rect -5105 -88 -5071 88
rect -5009 -88 -4975 88
rect -4913 -88 -4879 88
rect -4817 -88 -4783 88
rect -4721 -88 -4687 88
rect -4625 -88 -4591 88
rect -4529 -88 -4495 88
rect -4433 -88 -4399 88
rect -4337 -88 -4303 88
rect -4241 -88 -4207 88
rect -4145 -88 -4111 88
rect -4049 -88 -4015 88
rect -3953 -88 -3919 88
rect -3857 -88 -3823 88
rect -3761 -88 -3727 88
rect -3665 -88 -3631 88
rect -3569 -88 -3535 88
rect -3473 -88 -3439 88
rect -3377 -88 -3343 88
rect -3281 -88 -3247 88
rect -3185 -88 -3151 88
rect -3089 -88 -3055 88
rect -2993 -88 -2959 88
rect -2897 -88 -2863 88
rect -2801 -88 -2767 88
rect -2705 -88 -2671 88
rect -2609 -88 -2575 88
rect -2513 -88 -2479 88
rect -2417 -88 -2383 88
rect -2321 -88 -2287 88
rect -2225 -88 -2191 88
rect -2129 -88 -2095 88
rect -2033 -88 -1999 88
rect -1937 -88 -1903 88
rect -1841 -88 -1807 88
rect -1745 -88 -1711 88
rect -1649 -88 -1615 88
rect -1553 -88 -1519 88
rect -1457 -88 -1423 88
rect -1361 -88 -1327 88
rect -1265 -88 -1231 88
rect -1169 -88 -1135 88
rect -1073 -88 -1039 88
rect -977 -88 -943 88
rect -881 -88 -847 88
rect -785 -88 -751 88
rect -689 -88 -655 88
rect -593 -88 -559 88
rect -497 -88 -463 88
rect -401 -88 -367 88
rect -305 -88 -271 88
rect -209 -88 -175 88
rect -113 -88 -79 88
rect -17 -88 17 88
rect 79 -88 113 88
rect 175 -88 209 88
rect 271 -88 305 88
rect 367 -88 401 88
rect 463 -88 497 88
rect 559 -88 593 88
rect 655 -88 689 88
rect 751 -88 785 88
rect 847 -88 881 88
rect 943 -88 977 88
rect 1039 -88 1073 88
rect 1135 -88 1169 88
rect 1231 -88 1265 88
rect 1327 -88 1361 88
rect 1423 -88 1457 88
rect 1519 -88 1553 88
rect 1615 -88 1649 88
rect 1711 -88 1745 88
rect 1807 -88 1841 88
rect 1903 -88 1937 88
rect 1999 -88 2033 88
rect 2095 -88 2129 88
rect 2191 -88 2225 88
rect 2287 -88 2321 88
rect 2383 -88 2417 88
rect 2479 -88 2513 88
rect 2575 -88 2609 88
rect 2671 -88 2705 88
rect 2767 -88 2801 88
rect 2863 -88 2897 88
rect 2959 -88 2993 88
rect 3055 -88 3089 88
rect 3151 -88 3185 88
rect 3247 -88 3281 88
rect 3343 -88 3377 88
rect 3439 -88 3473 88
rect 3535 -88 3569 88
rect 3631 -88 3665 88
rect 3727 -88 3761 88
rect 3823 -88 3857 88
rect 3919 -88 3953 88
rect 4015 -88 4049 88
rect 4111 -88 4145 88
rect 4207 -88 4241 88
rect 4303 -88 4337 88
rect 4399 -88 4433 88
rect 4495 -88 4529 88
rect 4591 -88 4625 88
rect 4687 -88 4721 88
rect 4783 -88 4817 88
rect 4879 -88 4913 88
rect 4975 -88 5009 88
rect 5071 -88 5105 88
rect 5167 -88 5201 88
rect 5263 -88 5297 88
rect 5359 -88 5393 88
rect 5455 -88 5489 88
rect 5551 -88 5585 88
rect 5647 -88 5681 88
rect 5743 -88 5777 88
rect 5839 -88 5873 88
rect 5935 -88 5969 88
rect 6031 -88 6065 88
rect 6127 -88 6161 88
rect 6223 -88 6257 88
rect 6319 -88 6353 88
rect 6415 -88 6449 88
rect 6511 -88 6545 88
rect 6607 -88 6641 88
rect 6703 -88 6737 88
rect 6799 -88 6833 88
rect 6895 -88 6929 88
rect 6991 -88 7025 88
rect 7087 -88 7121 88
rect 7183 -88 7217 88
rect 7279 -88 7313 88
rect 7375 -88 7409 88
rect 7471 -88 7505 88
rect 7567 -88 7601 88
rect 7663 -88 7697 88
rect 7759 -88 7793 88
rect 7855 -88 7889 88
rect 7951 -88 7985 88
rect 8047 -88 8081 88
rect 8143 -88 8177 88
rect 8239 -88 8273 88
<< psubdiff >>
rect -8387 240 -8291 274
rect 8291 240 8387 274
rect -8387 178 -8353 240
rect 8353 178 8387 240
rect -8387 -240 -8353 -178
rect 8353 -240 8387 -178
rect -8387 -274 -8291 -240
rect 8291 -274 8387 -240
<< psubdiffcont >>
rect -8291 240 8291 274
rect -8387 -178 -8353 178
rect 8353 -178 8387 178
rect -8291 -274 8291 -240
<< poly >>
rect -8145 172 -8079 188
rect -8145 138 -8129 172
rect -8095 138 -8079 172
rect -8223 100 -8193 126
rect -8145 122 -8079 138
rect -7953 172 -7887 188
rect -7953 138 -7937 172
rect -7903 138 -7887 172
rect -8127 100 -8097 122
rect -8031 100 -8001 126
rect -7953 122 -7887 138
rect -7761 172 -7695 188
rect -7761 138 -7745 172
rect -7711 138 -7695 172
rect -7935 100 -7905 122
rect -7839 100 -7809 126
rect -7761 122 -7695 138
rect -7569 172 -7503 188
rect -7569 138 -7553 172
rect -7519 138 -7503 172
rect -7743 100 -7713 122
rect -7647 100 -7617 126
rect -7569 122 -7503 138
rect -7377 172 -7311 188
rect -7377 138 -7361 172
rect -7327 138 -7311 172
rect -7551 100 -7521 122
rect -7455 100 -7425 126
rect -7377 122 -7311 138
rect -7185 172 -7119 188
rect -7185 138 -7169 172
rect -7135 138 -7119 172
rect -7359 100 -7329 122
rect -7263 100 -7233 126
rect -7185 122 -7119 138
rect -6993 172 -6927 188
rect -6993 138 -6977 172
rect -6943 138 -6927 172
rect -7167 100 -7137 122
rect -7071 100 -7041 126
rect -6993 122 -6927 138
rect -6801 172 -6735 188
rect -6801 138 -6785 172
rect -6751 138 -6735 172
rect -6975 100 -6945 122
rect -6879 100 -6849 126
rect -6801 122 -6735 138
rect -6609 172 -6543 188
rect -6609 138 -6593 172
rect -6559 138 -6543 172
rect -6783 100 -6753 122
rect -6687 100 -6657 126
rect -6609 122 -6543 138
rect -6417 172 -6351 188
rect -6417 138 -6401 172
rect -6367 138 -6351 172
rect -6591 100 -6561 122
rect -6495 100 -6465 126
rect -6417 122 -6351 138
rect -6225 172 -6159 188
rect -6225 138 -6209 172
rect -6175 138 -6159 172
rect -6399 100 -6369 122
rect -6303 100 -6273 126
rect -6225 122 -6159 138
rect -6033 172 -5967 188
rect -6033 138 -6017 172
rect -5983 138 -5967 172
rect -6207 100 -6177 122
rect -6111 100 -6081 126
rect -6033 122 -5967 138
rect -5841 172 -5775 188
rect -5841 138 -5825 172
rect -5791 138 -5775 172
rect -6015 100 -5985 122
rect -5919 100 -5889 126
rect -5841 122 -5775 138
rect -5649 172 -5583 188
rect -5649 138 -5633 172
rect -5599 138 -5583 172
rect -5823 100 -5793 122
rect -5727 100 -5697 126
rect -5649 122 -5583 138
rect -5457 172 -5391 188
rect -5457 138 -5441 172
rect -5407 138 -5391 172
rect -5631 100 -5601 122
rect -5535 100 -5505 126
rect -5457 122 -5391 138
rect -5265 172 -5199 188
rect -5265 138 -5249 172
rect -5215 138 -5199 172
rect -5439 100 -5409 122
rect -5343 100 -5313 126
rect -5265 122 -5199 138
rect -5073 172 -5007 188
rect -5073 138 -5057 172
rect -5023 138 -5007 172
rect -5247 100 -5217 122
rect -5151 100 -5121 126
rect -5073 122 -5007 138
rect -4881 172 -4815 188
rect -4881 138 -4865 172
rect -4831 138 -4815 172
rect -5055 100 -5025 122
rect -4959 100 -4929 126
rect -4881 122 -4815 138
rect -4689 172 -4623 188
rect -4689 138 -4673 172
rect -4639 138 -4623 172
rect -4863 100 -4833 122
rect -4767 100 -4737 126
rect -4689 122 -4623 138
rect -4497 172 -4431 188
rect -4497 138 -4481 172
rect -4447 138 -4431 172
rect -4671 100 -4641 122
rect -4575 100 -4545 126
rect -4497 122 -4431 138
rect -4305 172 -4239 188
rect -4305 138 -4289 172
rect -4255 138 -4239 172
rect -4479 100 -4449 122
rect -4383 100 -4353 126
rect -4305 122 -4239 138
rect -4113 172 -4047 188
rect -4113 138 -4097 172
rect -4063 138 -4047 172
rect -4287 100 -4257 122
rect -4191 100 -4161 126
rect -4113 122 -4047 138
rect -3921 172 -3855 188
rect -3921 138 -3905 172
rect -3871 138 -3855 172
rect -4095 100 -4065 122
rect -3999 100 -3969 126
rect -3921 122 -3855 138
rect -3729 172 -3663 188
rect -3729 138 -3713 172
rect -3679 138 -3663 172
rect -3903 100 -3873 122
rect -3807 100 -3777 126
rect -3729 122 -3663 138
rect -3537 172 -3471 188
rect -3537 138 -3521 172
rect -3487 138 -3471 172
rect -3711 100 -3681 122
rect -3615 100 -3585 126
rect -3537 122 -3471 138
rect -3345 172 -3279 188
rect -3345 138 -3329 172
rect -3295 138 -3279 172
rect -3519 100 -3489 122
rect -3423 100 -3393 126
rect -3345 122 -3279 138
rect -3153 172 -3087 188
rect -3153 138 -3137 172
rect -3103 138 -3087 172
rect -3327 100 -3297 122
rect -3231 100 -3201 126
rect -3153 122 -3087 138
rect -2961 172 -2895 188
rect -2961 138 -2945 172
rect -2911 138 -2895 172
rect -3135 100 -3105 122
rect -3039 100 -3009 126
rect -2961 122 -2895 138
rect -2769 172 -2703 188
rect -2769 138 -2753 172
rect -2719 138 -2703 172
rect -2943 100 -2913 122
rect -2847 100 -2817 126
rect -2769 122 -2703 138
rect -2577 172 -2511 188
rect -2577 138 -2561 172
rect -2527 138 -2511 172
rect -2751 100 -2721 122
rect -2655 100 -2625 126
rect -2577 122 -2511 138
rect -2385 172 -2319 188
rect -2385 138 -2369 172
rect -2335 138 -2319 172
rect -2559 100 -2529 122
rect -2463 100 -2433 126
rect -2385 122 -2319 138
rect -2193 172 -2127 188
rect -2193 138 -2177 172
rect -2143 138 -2127 172
rect -2367 100 -2337 122
rect -2271 100 -2241 126
rect -2193 122 -2127 138
rect -2001 172 -1935 188
rect -2001 138 -1985 172
rect -1951 138 -1935 172
rect -2175 100 -2145 122
rect -2079 100 -2049 126
rect -2001 122 -1935 138
rect -1809 172 -1743 188
rect -1809 138 -1793 172
rect -1759 138 -1743 172
rect -1983 100 -1953 122
rect -1887 100 -1857 126
rect -1809 122 -1743 138
rect -1617 172 -1551 188
rect -1617 138 -1601 172
rect -1567 138 -1551 172
rect -1791 100 -1761 122
rect -1695 100 -1665 126
rect -1617 122 -1551 138
rect -1425 172 -1359 188
rect -1425 138 -1409 172
rect -1375 138 -1359 172
rect -1599 100 -1569 122
rect -1503 100 -1473 126
rect -1425 122 -1359 138
rect -1233 172 -1167 188
rect -1233 138 -1217 172
rect -1183 138 -1167 172
rect -1407 100 -1377 122
rect -1311 100 -1281 126
rect -1233 122 -1167 138
rect -1041 172 -975 188
rect -1041 138 -1025 172
rect -991 138 -975 172
rect -1215 100 -1185 122
rect -1119 100 -1089 126
rect -1041 122 -975 138
rect -849 172 -783 188
rect -849 138 -833 172
rect -799 138 -783 172
rect -1023 100 -993 122
rect -927 100 -897 126
rect -849 122 -783 138
rect -657 172 -591 188
rect -657 138 -641 172
rect -607 138 -591 172
rect -831 100 -801 122
rect -735 100 -705 126
rect -657 122 -591 138
rect -465 172 -399 188
rect -465 138 -449 172
rect -415 138 -399 172
rect -639 100 -609 122
rect -543 100 -513 126
rect -465 122 -399 138
rect -273 172 -207 188
rect -273 138 -257 172
rect -223 138 -207 172
rect -447 100 -417 122
rect -351 100 -321 126
rect -273 122 -207 138
rect -81 172 -15 188
rect -81 138 -65 172
rect -31 138 -15 172
rect -255 100 -225 122
rect -159 100 -129 126
rect -81 122 -15 138
rect 111 172 177 188
rect 111 138 127 172
rect 161 138 177 172
rect -63 100 -33 122
rect 33 100 63 126
rect 111 122 177 138
rect 303 172 369 188
rect 303 138 319 172
rect 353 138 369 172
rect 129 100 159 122
rect 225 100 255 126
rect 303 122 369 138
rect 495 172 561 188
rect 495 138 511 172
rect 545 138 561 172
rect 321 100 351 122
rect 417 100 447 126
rect 495 122 561 138
rect 687 172 753 188
rect 687 138 703 172
rect 737 138 753 172
rect 513 100 543 122
rect 609 100 639 126
rect 687 122 753 138
rect 879 172 945 188
rect 879 138 895 172
rect 929 138 945 172
rect 705 100 735 122
rect 801 100 831 126
rect 879 122 945 138
rect 1071 172 1137 188
rect 1071 138 1087 172
rect 1121 138 1137 172
rect 897 100 927 122
rect 993 100 1023 126
rect 1071 122 1137 138
rect 1263 172 1329 188
rect 1263 138 1279 172
rect 1313 138 1329 172
rect 1089 100 1119 122
rect 1185 100 1215 126
rect 1263 122 1329 138
rect 1455 172 1521 188
rect 1455 138 1471 172
rect 1505 138 1521 172
rect 1281 100 1311 122
rect 1377 100 1407 126
rect 1455 122 1521 138
rect 1647 172 1713 188
rect 1647 138 1663 172
rect 1697 138 1713 172
rect 1473 100 1503 122
rect 1569 100 1599 126
rect 1647 122 1713 138
rect 1839 172 1905 188
rect 1839 138 1855 172
rect 1889 138 1905 172
rect 1665 100 1695 122
rect 1761 100 1791 126
rect 1839 122 1905 138
rect 2031 172 2097 188
rect 2031 138 2047 172
rect 2081 138 2097 172
rect 1857 100 1887 122
rect 1953 100 1983 126
rect 2031 122 2097 138
rect 2223 172 2289 188
rect 2223 138 2239 172
rect 2273 138 2289 172
rect 2049 100 2079 122
rect 2145 100 2175 126
rect 2223 122 2289 138
rect 2415 172 2481 188
rect 2415 138 2431 172
rect 2465 138 2481 172
rect 2241 100 2271 122
rect 2337 100 2367 126
rect 2415 122 2481 138
rect 2607 172 2673 188
rect 2607 138 2623 172
rect 2657 138 2673 172
rect 2433 100 2463 122
rect 2529 100 2559 126
rect 2607 122 2673 138
rect 2799 172 2865 188
rect 2799 138 2815 172
rect 2849 138 2865 172
rect 2625 100 2655 122
rect 2721 100 2751 126
rect 2799 122 2865 138
rect 2991 172 3057 188
rect 2991 138 3007 172
rect 3041 138 3057 172
rect 2817 100 2847 122
rect 2913 100 2943 126
rect 2991 122 3057 138
rect 3183 172 3249 188
rect 3183 138 3199 172
rect 3233 138 3249 172
rect 3009 100 3039 122
rect 3105 100 3135 126
rect 3183 122 3249 138
rect 3375 172 3441 188
rect 3375 138 3391 172
rect 3425 138 3441 172
rect 3201 100 3231 122
rect 3297 100 3327 126
rect 3375 122 3441 138
rect 3567 172 3633 188
rect 3567 138 3583 172
rect 3617 138 3633 172
rect 3393 100 3423 122
rect 3489 100 3519 126
rect 3567 122 3633 138
rect 3759 172 3825 188
rect 3759 138 3775 172
rect 3809 138 3825 172
rect 3585 100 3615 122
rect 3681 100 3711 126
rect 3759 122 3825 138
rect 3951 172 4017 188
rect 3951 138 3967 172
rect 4001 138 4017 172
rect 3777 100 3807 122
rect 3873 100 3903 126
rect 3951 122 4017 138
rect 4143 172 4209 188
rect 4143 138 4159 172
rect 4193 138 4209 172
rect 3969 100 3999 122
rect 4065 100 4095 126
rect 4143 122 4209 138
rect 4335 172 4401 188
rect 4335 138 4351 172
rect 4385 138 4401 172
rect 4161 100 4191 122
rect 4257 100 4287 126
rect 4335 122 4401 138
rect 4527 172 4593 188
rect 4527 138 4543 172
rect 4577 138 4593 172
rect 4353 100 4383 122
rect 4449 100 4479 126
rect 4527 122 4593 138
rect 4719 172 4785 188
rect 4719 138 4735 172
rect 4769 138 4785 172
rect 4545 100 4575 122
rect 4641 100 4671 126
rect 4719 122 4785 138
rect 4911 172 4977 188
rect 4911 138 4927 172
rect 4961 138 4977 172
rect 4737 100 4767 122
rect 4833 100 4863 126
rect 4911 122 4977 138
rect 5103 172 5169 188
rect 5103 138 5119 172
rect 5153 138 5169 172
rect 4929 100 4959 122
rect 5025 100 5055 126
rect 5103 122 5169 138
rect 5295 172 5361 188
rect 5295 138 5311 172
rect 5345 138 5361 172
rect 5121 100 5151 122
rect 5217 100 5247 126
rect 5295 122 5361 138
rect 5487 172 5553 188
rect 5487 138 5503 172
rect 5537 138 5553 172
rect 5313 100 5343 122
rect 5409 100 5439 126
rect 5487 122 5553 138
rect 5679 172 5745 188
rect 5679 138 5695 172
rect 5729 138 5745 172
rect 5505 100 5535 122
rect 5601 100 5631 126
rect 5679 122 5745 138
rect 5871 172 5937 188
rect 5871 138 5887 172
rect 5921 138 5937 172
rect 5697 100 5727 122
rect 5793 100 5823 126
rect 5871 122 5937 138
rect 6063 172 6129 188
rect 6063 138 6079 172
rect 6113 138 6129 172
rect 5889 100 5919 122
rect 5985 100 6015 126
rect 6063 122 6129 138
rect 6255 172 6321 188
rect 6255 138 6271 172
rect 6305 138 6321 172
rect 6081 100 6111 122
rect 6177 100 6207 126
rect 6255 122 6321 138
rect 6447 172 6513 188
rect 6447 138 6463 172
rect 6497 138 6513 172
rect 6273 100 6303 122
rect 6369 100 6399 126
rect 6447 122 6513 138
rect 6639 172 6705 188
rect 6639 138 6655 172
rect 6689 138 6705 172
rect 6465 100 6495 122
rect 6561 100 6591 126
rect 6639 122 6705 138
rect 6831 172 6897 188
rect 6831 138 6847 172
rect 6881 138 6897 172
rect 6657 100 6687 122
rect 6753 100 6783 126
rect 6831 122 6897 138
rect 7023 172 7089 188
rect 7023 138 7039 172
rect 7073 138 7089 172
rect 6849 100 6879 122
rect 6945 100 6975 126
rect 7023 122 7089 138
rect 7215 172 7281 188
rect 7215 138 7231 172
rect 7265 138 7281 172
rect 7041 100 7071 122
rect 7137 100 7167 126
rect 7215 122 7281 138
rect 7407 172 7473 188
rect 7407 138 7423 172
rect 7457 138 7473 172
rect 7233 100 7263 122
rect 7329 100 7359 126
rect 7407 122 7473 138
rect 7599 172 7665 188
rect 7599 138 7615 172
rect 7649 138 7665 172
rect 7425 100 7455 122
rect 7521 100 7551 126
rect 7599 122 7665 138
rect 7791 172 7857 188
rect 7791 138 7807 172
rect 7841 138 7857 172
rect 7617 100 7647 122
rect 7713 100 7743 126
rect 7791 122 7857 138
rect 7983 172 8049 188
rect 7983 138 7999 172
rect 8033 138 8049 172
rect 7809 100 7839 122
rect 7905 100 7935 126
rect 7983 122 8049 138
rect 8175 172 8241 188
rect 8175 138 8191 172
rect 8225 138 8241 172
rect 8001 100 8031 122
rect 8097 100 8127 126
rect 8175 122 8241 138
rect 8193 100 8223 122
rect -8223 -122 -8193 -100
rect -8241 -138 -8175 -122
rect -8127 -126 -8097 -100
rect -8031 -122 -8001 -100
rect -8241 -172 -8225 -138
rect -8191 -172 -8175 -138
rect -8241 -188 -8175 -172
rect -8049 -138 -7983 -122
rect -7935 -126 -7905 -100
rect -7839 -122 -7809 -100
rect -8049 -172 -8033 -138
rect -7999 -172 -7983 -138
rect -8049 -188 -7983 -172
rect -7857 -138 -7791 -122
rect -7743 -126 -7713 -100
rect -7647 -122 -7617 -100
rect -7857 -172 -7841 -138
rect -7807 -172 -7791 -138
rect -7857 -188 -7791 -172
rect -7665 -138 -7599 -122
rect -7551 -126 -7521 -100
rect -7455 -122 -7425 -100
rect -7665 -172 -7649 -138
rect -7615 -172 -7599 -138
rect -7665 -188 -7599 -172
rect -7473 -138 -7407 -122
rect -7359 -126 -7329 -100
rect -7263 -122 -7233 -100
rect -7473 -172 -7457 -138
rect -7423 -172 -7407 -138
rect -7473 -188 -7407 -172
rect -7281 -138 -7215 -122
rect -7167 -126 -7137 -100
rect -7071 -122 -7041 -100
rect -7281 -172 -7265 -138
rect -7231 -172 -7215 -138
rect -7281 -188 -7215 -172
rect -7089 -138 -7023 -122
rect -6975 -126 -6945 -100
rect -6879 -122 -6849 -100
rect -7089 -172 -7073 -138
rect -7039 -172 -7023 -138
rect -7089 -188 -7023 -172
rect -6897 -138 -6831 -122
rect -6783 -126 -6753 -100
rect -6687 -122 -6657 -100
rect -6897 -172 -6881 -138
rect -6847 -172 -6831 -138
rect -6897 -188 -6831 -172
rect -6705 -138 -6639 -122
rect -6591 -126 -6561 -100
rect -6495 -122 -6465 -100
rect -6705 -172 -6689 -138
rect -6655 -172 -6639 -138
rect -6705 -188 -6639 -172
rect -6513 -138 -6447 -122
rect -6399 -126 -6369 -100
rect -6303 -122 -6273 -100
rect -6513 -172 -6497 -138
rect -6463 -172 -6447 -138
rect -6513 -188 -6447 -172
rect -6321 -138 -6255 -122
rect -6207 -126 -6177 -100
rect -6111 -122 -6081 -100
rect -6321 -172 -6305 -138
rect -6271 -172 -6255 -138
rect -6321 -188 -6255 -172
rect -6129 -138 -6063 -122
rect -6015 -126 -5985 -100
rect -5919 -122 -5889 -100
rect -6129 -172 -6113 -138
rect -6079 -172 -6063 -138
rect -6129 -188 -6063 -172
rect -5937 -138 -5871 -122
rect -5823 -126 -5793 -100
rect -5727 -122 -5697 -100
rect -5937 -172 -5921 -138
rect -5887 -172 -5871 -138
rect -5937 -188 -5871 -172
rect -5745 -138 -5679 -122
rect -5631 -126 -5601 -100
rect -5535 -122 -5505 -100
rect -5745 -172 -5729 -138
rect -5695 -172 -5679 -138
rect -5745 -188 -5679 -172
rect -5553 -138 -5487 -122
rect -5439 -126 -5409 -100
rect -5343 -122 -5313 -100
rect -5553 -172 -5537 -138
rect -5503 -172 -5487 -138
rect -5553 -188 -5487 -172
rect -5361 -138 -5295 -122
rect -5247 -126 -5217 -100
rect -5151 -122 -5121 -100
rect -5361 -172 -5345 -138
rect -5311 -172 -5295 -138
rect -5361 -188 -5295 -172
rect -5169 -138 -5103 -122
rect -5055 -126 -5025 -100
rect -4959 -122 -4929 -100
rect -5169 -172 -5153 -138
rect -5119 -172 -5103 -138
rect -5169 -188 -5103 -172
rect -4977 -138 -4911 -122
rect -4863 -126 -4833 -100
rect -4767 -122 -4737 -100
rect -4977 -172 -4961 -138
rect -4927 -172 -4911 -138
rect -4977 -188 -4911 -172
rect -4785 -138 -4719 -122
rect -4671 -126 -4641 -100
rect -4575 -122 -4545 -100
rect -4785 -172 -4769 -138
rect -4735 -172 -4719 -138
rect -4785 -188 -4719 -172
rect -4593 -138 -4527 -122
rect -4479 -126 -4449 -100
rect -4383 -122 -4353 -100
rect -4593 -172 -4577 -138
rect -4543 -172 -4527 -138
rect -4593 -188 -4527 -172
rect -4401 -138 -4335 -122
rect -4287 -126 -4257 -100
rect -4191 -122 -4161 -100
rect -4401 -172 -4385 -138
rect -4351 -172 -4335 -138
rect -4401 -188 -4335 -172
rect -4209 -138 -4143 -122
rect -4095 -126 -4065 -100
rect -3999 -122 -3969 -100
rect -4209 -172 -4193 -138
rect -4159 -172 -4143 -138
rect -4209 -188 -4143 -172
rect -4017 -138 -3951 -122
rect -3903 -126 -3873 -100
rect -3807 -122 -3777 -100
rect -4017 -172 -4001 -138
rect -3967 -172 -3951 -138
rect -4017 -188 -3951 -172
rect -3825 -138 -3759 -122
rect -3711 -126 -3681 -100
rect -3615 -122 -3585 -100
rect -3825 -172 -3809 -138
rect -3775 -172 -3759 -138
rect -3825 -188 -3759 -172
rect -3633 -138 -3567 -122
rect -3519 -126 -3489 -100
rect -3423 -122 -3393 -100
rect -3633 -172 -3617 -138
rect -3583 -172 -3567 -138
rect -3633 -188 -3567 -172
rect -3441 -138 -3375 -122
rect -3327 -126 -3297 -100
rect -3231 -122 -3201 -100
rect -3441 -172 -3425 -138
rect -3391 -172 -3375 -138
rect -3441 -188 -3375 -172
rect -3249 -138 -3183 -122
rect -3135 -126 -3105 -100
rect -3039 -122 -3009 -100
rect -3249 -172 -3233 -138
rect -3199 -172 -3183 -138
rect -3249 -188 -3183 -172
rect -3057 -138 -2991 -122
rect -2943 -126 -2913 -100
rect -2847 -122 -2817 -100
rect -3057 -172 -3041 -138
rect -3007 -172 -2991 -138
rect -3057 -188 -2991 -172
rect -2865 -138 -2799 -122
rect -2751 -126 -2721 -100
rect -2655 -122 -2625 -100
rect -2865 -172 -2849 -138
rect -2815 -172 -2799 -138
rect -2865 -188 -2799 -172
rect -2673 -138 -2607 -122
rect -2559 -126 -2529 -100
rect -2463 -122 -2433 -100
rect -2673 -172 -2657 -138
rect -2623 -172 -2607 -138
rect -2673 -188 -2607 -172
rect -2481 -138 -2415 -122
rect -2367 -126 -2337 -100
rect -2271 -122 -2241 -100
rect -2481 -172 -2465 -138
rect -2431 -172 -2415 -138
rect -2481 -188 -2415 -172
rect -2289 -138 -2223 -122
rect -2175 -126 -2145 -100
rect -2079 -122 -2049 -100
rect -2289 -172 -2273 -138
rect -2239 -172 -2223 -138
rect -2289 -188 -2223 -172
rect -2097 -138 -2031 -122
rect -1983 -126 -1953 -100
rect -1887 -122 -1857 -100
rect -2097 -172 -2081 -138
rect -2047 -172 -2031 -138
rect -2097 -188 -2031 -172
rect -1905 -138 -1839 -122
rect -1791 -126 -1761 -100
rect -1695 -122 -1665 -100
rect -1905 -172 -1889 -138
rect -1855 -172 -1839 -138
rect -1905 -188 -1839 -172
rect -1713 -138 -1647 -122
rect -1599 -126 -1569 -100
rect -1503 -122 -1473 -100
rect -1713 -172 -1697 -138
rect -1663 -172 -1647 -138
rect -1713 -188 -1647 -172
rect -1521 -138 -1455 -122
rect -1407 -126 -1377 -100
rect -1311 -122 -1281 -100
rect -1521 -172 -1505 -138
rect -1471 -172 -1455 -138
rect -1521 -188 -1455 -172
rect -1329 -138 -1263 -122
rect -1215 -126 -1185 -100
rect -1119 -122 -1089 -100
rect -1329 -172 -1313 -138
rect -1279 -172 -1263 -138
rect -1329 -188 -1263 -172
rect -1137 -138 -1071 -122
rect -1023 -126 -993 -100
rect -927 -122 -897 -100
rect -1137 -172 -1121 -138
rect -1087 -172 -1071 -138
rect -1137 -188 -1071 -172
rect -945 -138 -879 -122
rect -831 -126 -801 -100
rect -735 -122 -705 -100
rect -945 -172 -929 -138
rect -895 -172 -879 -138
rect -945 -188 -879 -172
rect -753 -138 -687 -122
rect -639 -126 -609 -100
rect -543 -122 -513 -100
rect -753 -172 -737 -138
rect -703 -172 -687 -138
rect -753 -188 -687 -172
rect -561 -138 -495 -122
rect -447 -126 -417 -100
rect -351 -122 -321 -100
rect -561 -172 -545 -138
rect -511 -172 -495 -138
rect -561 -188 -495 -172
rect -369 -138 -303 -122
rect -255 -126 -225 -100
rect -159 -122 -129 -100
rect -369 -172 -353 -138
rect -319 -172 -303 -138
rect -369 -188 -303 -172
rect -177 -138 -111 -122
rect -63 -126 -33 -100
rect 33 -122 63 -100
rect -177 -172 -161 -138
rect -127 -172 -111 -138
rect -177 -188 -111 -172
rect 15 -138 81 -122
rect 129 -126 159 -100
rect 225 -122 255 -100
rect 15 -172 31 -138
rect 65 -172 81 -138
rect 15 -188 81 -172
rect 207 -138 273 -122
rect 321 -126 351 -100
rect 417 -122 447 -100
rect 207 -172 223 -138
rect 257 -172 273 -138
rect 207 -188 273 -172
rect 399 -138 465 -122
rect 513 -126 543 -100
rect 609 -122 639 -100
rect 399 -172 415 -138
rect 449 -172 465 -138
rect 399 -188 465 -172
rect 591 -138 657 -122
rect 705 -126 735 -100
rect 801 -122 831 -100
rect 591 -172 607 -138
rect 641 -172 657 -138
rect 591 -188 657 -172
rect 783 -138 849 -122
rect 897 -126 927 -100
rect 993 -122 1023 -100
rect 783 -172 799 -138
rect 833 -172 849 -138
rect 783 -188 849 -172
rect 975 -138 1041 -122
rect 1089 -126 1119 -100
rect 1185 -122 1215 -100
rect 975 -172 991 -138
rect 1025 -172 1041 -138
rect 975 -188 1041 -172
rect 1167 -138 1233 -122
rect 1281 -126 1311 -100
rect 1377 -122 1407 -100
rect 1167 -172 1183 -138
rect 1217 -172 1233 -138
rect 1167 -188 1233 -172
rect 1359 -138 1425 -122
rect 1473 -126 1503 -100
rect 1569 -122 1599 -100
rect 1359 -172 1375 -138
rect 1409 -172 1425 -138
rect 1359 -188 1425 -172
rect 1551 -138 1617 -122
rect 1665 -126 1695 -100
rect 1761 -122 1791 -100
rect 1551 -172 1567 -138
rect 1601 -172 1617 -138
rect 1551 -188 1617 -172
rect 1743 -138 1809 -122
rect 1857 -126 1887 -100
rect 1953 -122 1983 -100
rect 1743 -172 1759 -138
rect 1793 -172 1809 -138
rect 1743 -188 1809 -172
rect 1935 -138 2001 -122
rect 2049 -126 2079 -100
rect 2145 -122 2175 -100
rect 1935 -172 1951 -138
rect 1985 -172 2001 -138
rect 1935 -188 2001 -172
rect 2127 -138 2193 -122
rect 2241 -126 2271 -100
rect 2337 -122 2367 -100
rect 2127 -172 2143 -138
rect 2177 -172 2193 -138
rect 2127 -188 2193 -172
rect 2319 -138 2385 -122
rect 2433 -126 2463 -100
rect 2529 -122 2559 -100
rect 2319 -172 2335 -138
rect 2369 -172 2385 -138
rect 2319 -188 2385 -172
rect 2511 -138 2577 -122
rect 2625 -126 2655 -100
rect 2721 -122 2751 -100
rect 2511 -172 2527 -138
rect 2561 -172 2577 -138
rect 2511 -188 2577 -172
rect 2703 -138 2769 -122
rect 2817 -126 2847 -100
rect 2913 -122 2943 -100
rect 2703 -172 2719 -138
rect 2753 -172 2769 -138
rect 2703 -188 2769 -172
rect 2895 -138 2961 -122
rect 3009 -126 3039 -100
rect 3105 -122 3135 -100
rect 2895 -172 2911 -138
rect 2945 -172 2961 -138
rect 2895 -188 2961 -172
rect 3087 -138 3153 -122
rect 3201 -126 3231 -100
rect 3297 -122 3327 -100
rect 3087 -172 3103 -138
rect 3137 -172 3153 -138
rect 3087 -188 3153 -172
rect 3279 -138 3345 -122
rect 3393 -126 3423 -100
rect 3489 -122 3519 -100
rect 3279 -172 3295 -138
rect 3329 -172 3345 -138
rect 3279 -188 3345 -172
rect 3471 -138 3537 -122
rect 3585 -126 3615 -100
rect 3681 -122 3711 -100
rect 3471 -172 3487 -138
rect 3521 -172 3537 -138
rect 3471 -188 3537 -172
rect 3663 -138 3729 -122
rect 3777 -126 3807 -100
rect 3873 -122 3903 -100
rect 3663 -172 3679 -138
rect 3713 -172 3729 -138
rect 3663 -188 3729 -172
rect 3855 -138 3921 -122
rect 3969 -126 3999 -100
rect 4065 -122 4095 -100
rect 3855 -172 3871 -138
rect 3905 -172 3921 -138
rect 3855 -188 3921 -172
rect 4047 -138 4113 -122
rect 4161 -126 4191 -100
rect 4257 -122 4287 -100
rect 4047 -172 4063 -138
rect 4097 -172 4113 -138
rect 4047 -188 4113 -172
rect 4239 -138 4305 -122
rect 4353 -126 4383 -100
rect 4449 -122 4479 -100
rect 4239 -172 4255 -138
rect 4289 -172 4305 -138
rect 4239 -188 4305 -172
rect 4431 -138 4497 -122
rect 4545 -126 4575 -100
rect 4641 -122 4671 -100
rect 4431 -172 4447 -138
rect 4481 -172 4497 -138
rect 4431 -188 4497 -172
rect 4623 -138 4689 -122
rect 4737 -126 4767 -100
rect 4833 -122 4863 -100
rect 4623 -172 4639 -138
rect 4673 -172 4689 -138
rect 4623 -188 4689 -172
rect 4815 -138 4881 -122
rect 4929 -126 4959 -100
rect 5025 -122 5055 -100
rect 4815 -172 4831 -138
rect 4865 -172 4881 -138
rect 4815 -188 4881 -172
rect 5007 -138 5073 -122
rect 5121 -126 5151 -100
rect 5217 -122 5247 -100
rect 5007 -172 5023 -138
rect 5057 -172 5073 -138
rect 5007 -188 5073 -172
rect 5199 -138 5265 -122
rect 5313 -126 5343 -100
rect 5409 -122 5439 -100
rect 5199 -172 5215 -138
rect 5249 -172 5265 -138
rect 5199 -188 5265 -172
rect 5391 -138 5457 -122
rect 5505 -126 5535 -100
rect 5601 -122 5631 -100
rect 5391 -172 5407 -138
rect 5441 -172 5457 -138
rect 5391 -188 5457 -172
rect 5583 -138 5649 -122
rect 5697 -126 5727 -100
rect 5793 -122 5823 -100
rect 5583 -172 5599 -138
rect 5633 -172 5649 -138
rect 5583 -188 5649 -172
rect 5775 -138 5841 -122
rect 5889 -126 5919 -100
rect 5985 -122 6015 -100
rect 5775 -172 5791 -138
rect 5825 -172 5841 -138
rect 5775 -188 5841 -172
rect 5967 -138 6033 -122
rect 6081 -126 6111 -100
rect 6177 -122 6207 -100
rect 5967 -172 5983 -138
rect 6017 -172 6033 -138
rect 5967 -188 6033 -172
rect 6159 -138 6225 -122
rect 6273 -126 6303 -100
rect 6369 -122 6399 -100
rect 6159 -172 6175 -138
rect 6209 -172 6225 -138
rect 6159 -188 6225 -172
rect 6351 -138 6417 -122
rect 6465 -126 6495 -100
rect 6561 -122 6591 -100
rect 6351 -172 6367 -138
rect 6401 -172 6417 -138
rect 6351 -188 6417 -172
rect 6543 -138 6609 -122
rect 6657 -126 6687 -100
rect 6753 -122 6783 -100
rect 6543 -172 6559 -138
rect 6593 -172 6609 -138
rect 6543 -188 6609 -172
rect 6735 -138 6801 -122
rect 6849 -126 6879 -100
rect 6945 -122 6975 -100
rect 6735 -172 6751 -138
rect 6785 -172 6801 -138
rect 6735 -188 6801 -172
rect 6927 -138 6993 -122
rect 7041 -126 7071 -100
rect 7137 -122 7167 -100
rect 6927 -172 6943 -138
rect 6977 -172 6993 -138
rect 6927 -188 6993 -172
rect 7119 -138 7185 -122
rect 7233 -126 7263 -100
rect 7329 -122 7359 -100
rect 7119 -172 7135 -138
rect 7169 -172 7185 -138
rect 7119 -188 7185 -172
rect 7311 -138 7377 -122
rect 7425 -126 7455 -100
rect 7521 -122 7551 -100
rect 7311 -172 7327 -138
rect 7361 -172 7377 -138
rect 7311 -188 7377 -172
rect 7503 -138 7569 -122
rect 7617 -126 7647 -100
rect 7713 -122 7743 -100
rect 7503 -172 7519 -138
rect 7553 -172 7569 -138
rect 7503 -188 7569 -172
rect 7695 -138 7761 -122
rect 7809 -126 7839 -100
rect 7905 -122 7935 -100
rect 7695 -172 7711 -138
rect 7745 -172 7761 -138
rect 7695 -188 7761 -172
rect 7887 -138 7953 -122
rect 8001 -126 8031 -100
rect 8097 -122 8127 -100
rect 7887 -172 7903 -138
rect 7937 -172 7953 -138
rect 7887 -188 7953 -172
rect 8079 -138 8145 -122
rect 8193 -126 8223 -100
rect 8079 -172 8095 -138
rect 8129 -172 8145 -138
rect 8079 -188 8145 -172
<< polycont >>
rect -8129 138 -8095 172
rect -7937 138 -7903 172
rect -7745 138 -7711 172
rect -7553 138 -7519 172
rect -7361 138 -7327 172
rect -7169 138 -7135 172
rect -6977 138 -6943 172
rect -6785 138 -6751 172
rect -6593 138 -6559 172
rect -6401 138 -6367 172
rect -6209 138 -6175 172
rect -6017 138 -5983 172
rect -5825 138 -5791 172
rect -5633 138 -5599 172
rect -5441 138 -5407 172
rect -5249 138 -5215 172
rect -5057 138 -5023 172
rect -4865 138 -4831 172
rect -4673 138 -4639 172
rect -4481 138 -4447 172
rect -4289 138 -4255 172
rect -4097 138 -4063 172
rect -3905 138 -3871 172
rect -3713 138 -3679 172
rect -3521 138 -3487 172
rect -3329 138 -3295 172
rect -3137 138 -3103 172
rect -2945 138 -2911 172
rect -2753 138 -2719 172
rect -2561 138 -2527 172
rect -2369 138 -2335 172
rect -2177 138 -2143 172
rect -1985 138 -1951 172
rect -1793 138 -1759 172
rect -1601 138 -1567 172
rect -1409 138 -1375 172
rect -1217 138 -1183 172
rect -1025 138 -991 172
rect -833 138 -799 172
rect -641 138 -607 172
rect -449 138 -415 172
rect -257 138 -223 172
rect -65 138 -31 172
rect 127 138 161 172
rect 319 138 353 172
rect 511 138 545 172
rect 703 138 737 172
rect 895 138 929 172
rect 1087 138 1121 172
rect 1279 138 1313 172
rect 1471 138 1505 172
rect 1663 138 1697 172
rect 1855 138 1889 172
rect 2047 138 2081 172
rect 2239 138 2273 172
rect 2431 138 2465 172
rect 2623 138 2657 172
rect 2815 138 2849 172
rect 3007 138 3041 172
rect 3199 138 3233 172
rect 3391 138 3425 172
rect 3583 138 3617 172
rect 3775 138 3809 172
rect 3967 138 4001 172
rect 4159 138 4193 172
rect 4351 138 4385 172
rect 4543 138 4577 172
rect 4735 138 4769 172
rect 4927 138 4961 172
rect 5119 138 5153 172
rect 5311 138 5345 172
rect 5503 138 5537 172
rect 5695 138 5729 172
rect 5887 138 5921 172
rect 6079 138 6113 172
rect 6271 138 6305 172
rect 6463 138 6497 172
rect 6655 138 6689 172
rect 6847 138 6881 172
rect 7039 138 7073 172
rect 7231 138 7265 172
rect 7423 138 7457 172
rect 7615 138 7649 172
rect 7807 138 7841 172
rect 7999 138 8033 172
rect 8191 138 8225 172
rect -8225 -172 -8191 -138
rect -8033 -172 -7999 -138
rect -7841 -172 -7807 -138
rect -7649 -172 -7615 -138
rect -7457 -172 -7423 -138
rect -7265 -172 -7231 -138
rect -7073 -172 -7039 -138
rect -6881 -172 -6847 -138
rect -6689 -172 -6655 -138
rect -6497 -172 -6463 -138
rect -6305 -172 -6271 -138
rect -6113 -172 -6079 -138
rect -5921 -172 -5887 -138
rect -5729 -172 -5695 -138
rect -5537 -172 -5503 -138
rect -5345 -172 -5311 -138
rect -5153 -172 -5119 -138
rect -4961 -172 -4927 -138
rect -4769 -172 -4735 -138
rect -4577 -172 -4543 -138
rect -4385 -172 -4351 -138
rect -4193 -172 -4159 -138
rect -4001 -172 -3967 -138
rect -3809 -172 -3775 -138
rect -3617 -172 -3583 -138
rect -3425 -172 -3391 -138
rect -3233 -172 -3199 -138
rect -3041 -172 -3007 -138
rect -2849 -172 -2815 -138
rect -2657 -172 -2623 -138
rect -2465 -172 -2431 -138
rect -2273 -172 -2239 -138
rect -2081 -172 -2047 -138
rect -1889 -172 -1855 -138
rect -1697 -172 -1663 -138
rect -1505 -172 -1471 -138
rect -1313 -172 -1279 -138
rect -1121 -172 -1087 -138
rect -929 -172 -895 -138
rect -737 -172 -703 -138
rect -545 -172 -511 -138
rect -353 -172 -319 -138
rect -161 -172 -127 -138
rect 31 -172 65 -138
rect 223 -172 257 -138
rect 415 -172 449 -138
rect 607 -172 641 -138
rect 799 -172 833 -138
rect 991 -172 1025 -138
rect 1183 -172 1217 -138
rect 1375 -172 1409 -138
rect 1567 -172 1601 -138
rect 1759 -172 1793 -138
rect 1951 -172 1985 -138
rect 2143 -172 2177 -138
rect 2335 -172 2369 -138
rect 2527 -172 2561 -138
rect 2719 -172 2753 -138
rect 2911 -172 2945 -138
rect 3103 -172 3137 -138
rect 3295 -172 3329 -138
rect 3487 -172 3521 -138
rect 3679 -172 3713 -138
rect 3871 -172 3905 -138
rect 4063 -172 4097 -138
rect 4255 -172 4289 -138
rect 4447 -172 4481 -138
rect 4639 -172 4673 -138
rect 4831 -172 4865 -138
rect 5023 -172 5057 -138
rect 5215 -172 5249 -138
rect 5407 -172 5441 -138
rect 5599 -172 5633 -138
rect 5791 -172 5825 -138
rect 5983 -172 6017 -138
rect 6175 -172 6209 -138
rect 6367 -172 6401 -138
rect 6559 -172 6593 -138
rect 6751 -172 6785 -138
rect 6943 -172 6977 -138
rect 7135 -172 7169 -138
rect 7327 -172 7361 -138
rect 7519 -172 7553 -138
rect 7711 -172 7745 -138
rect 7903 -172 7937 -138
rect 8095 -172 8129 -138
<< locali >>
rect -8387 240 -8291 274
rect 8291 240 8387 274
rect -8387 178 -8353 240
rect 8353 178 8387 240
rect -8145 138 -8129 172
rect -8095 138 -8079 172
rect -7953 138 -7937 172
rect -7903 138 -7887 172
rect -7761 138 -7745 172
rect -7711 138 -7695 172
rect -7569 138 -7553 172
rect -7519 138 -7503 172
rect -7377 138 -7361 172
rect -7327 138 -7311 172
rect -7185 138 -7169 172
rect -7135 138 -7119 172
rect -6993 138 -6977 172
rect -6943 138 -6927 172
rect -6801 138 -6785 172
rect -6751 138 -6735 172
rect -6609 138 -6593 172
rect -6559 138 -6543 172
rect -6417 138 -6401 172
rect -6367 138 -6351 172
rect -6225 138 -6209 172
rect -6175 138 -6159 172
rect -6033 138 -6017 172
rect -5983 138 -5967 172
rect -5841 138 -5825 172
rect -5791 138 -5775 172
rect -5649 138 -5633 172
rect -5599 138 -5583 172
rect -5457 138 -5441 172
rect -5407 138 -5391 172
rect -5265 138 -5249 172
rect -5215 138 -5199 172
rect -5073 138 -5057 172
rect -5023 138 -5007 172
rect -4881 138 -4865 172
rect -4831 138 -4815 172
rect -4689 138 -4673 172
rect -4639 138 -4623 172
rect -4497 138 -4481 172
rect -4447 138 -4431 172
rect -4305 138 -4289 172
rect -4255 138 -4239 172
rect -4113 138 -4097 172
rect -4063 138 -4047 172
rect -3921 138 -3905 172
rect -3871 138 -3855 172
rect -3729 138 -3713 172
rect -3679 138 -3663 172
rect -3537 138 -3521 172
rect -3487 138 -3471 172
rect -3345 138 -3329 172
rect -3295 138 -3279 172
rect -3153 138 -3137 172
rect -3103 138 -3087 172
rect -2961 138 -2945 172
rect -2911 138 -2895 172
rect -2769 138 -2753 172
rect -2719 138 -2703 172
rect -2577 138 -2561 172
rect -2527 138 -2511 172
rect -2385 138 -2369 172
rect -2335 138 -2319 172
rect -2193 138 -2177 172
rect -2143 138 -2127 172
rect -2001 138 -1985 172
rect -1951 138 -1935 172
rect -1809 138 -1793 172
rect -1759 138 -1743 172
rect -1617 138 -1601 172
rect -1567 138 -1551 172
rect -1425 138 -1409 172
rect -1375 138 -1359 172
rect -1233 138 -1217 172
rect -1183 138 -1167 172
rect -1041 138 -1025 172
rect -991 138 -975 172
rect -849 138 -833 172
rect -799 138 -783 172
rect -657 138 -641 172
rect -607 138 -591 172
rect -465 138 -449 172
rect -415 138 -399 172
rect -273 138 -257 172
rect -223 138 -207 172
rect -81 138 -65 172
rect -31 138 -15 172
rect 111 138 127 172
rect 161 138 177 172
rect 303 138 319 172
rect 353 138 369 172
rect 495 138 511 172
rect 545 138 561 172
rect 687 138 703 172
rect 737 138 753 172
rect 879 138 895 172
rect 929 138 945 172
rect 1071 138 1087 172
rect 1121 138 1137 172
rect 1263 138 1279 172
rect 1313 138 1329 172
rect 1455 138 1471 172
rect 1505 138 1521 172
rect 1647 138 1663 172
rect 1697 138 1713 172
rect 1839 138 1855 172
rect 1889 138 1905 172
rect 2031 138 2047 172
rect 2081 138 2097 172
rect 2223 138 2239 172
rect 2273 138 2289 172
rect 2415 138 2431 172
rect 2465 138 2481 172
rect 2607 138 2623 172
rect 2657 138 2673 172
rect 2799 138 2815 172
rect 2849 138 2865 172
rect 2991 138 3007 172
rect 3041 138 3057 172
rect 3183 138 3199 172
rect 3233 138 3249 172
rect 3375 138 3391 172
rect 3425 138 3441 172
rect 3567 138 3583 172
rect 3617 138 3633 172
rect 3759 138 3775 172
rect 3809 138 3825 172
rect 3951 138 3967 172
rect 4001 138 4017 172
rect 4143 138 4159 172
rect 4193 138 4209 172
rect 4335 138 4351 172
rect 4385 138 4401 172
rect 4527 138 4543 172
rect 4577 138 4593 172
rect 4719 138 4735 172
rect 4769 138 4785 172
rect 4911 138 4927 172
rect 4961 138 4977 172
rect 5103 138 5119 172
rect 5153 138 5169 172
rect 5295 138 5311 172
rect 5345 138 5361 172
rect 5487 138 5503 172
rect 5537 138 5553 172
rect 5679 138 5695 172
rect 5729 138 5745 172
rect 5871 138 5887 172
rect 5921 138 5937 172
rect 6063 138 6079 172
rect 6113 138 6129 172
rect 6255 138 6271 172
rect 6305 138 6321 172
rect 6447 138 6463 172
rect 6497 138 6513 172
rect 6639 138 6655 172
rect 6689 138 6705 172
rect 6831 138 6847 172
rect 6881 138 6897 172
rect 7023 138 7039 172
rect 7073 138 7089 172
rect 7215 138 7231 172
rect 7265 138 7281 172
rect 7407 138 7423 172
rect 7457 138 7473 172
rect 7599 138 7615 172
rect 7649 138 7665 172
rect 7791 138 7807 172
rect 7841 138 7857 172
rect 7983 138 7999 172
rect 8033 138 8049 172
rect 8175 138 8191 172
rect 8225 138 8241 172
rect -8273 88 -8239 104
rect -8273 -104 -8239 -88
rect -8177 88 -8143 104
rect -8177 -104 -8143 -88
rect -8081 88 -8047 104
rect -8081 -104 -8047 -88
rect -7985 88 -7951 104
rect -7985 -104 -7951 -88
rect -7889 88 -7855 104
rect -7889 -104 -7855 -88
rect -7793 88 -7759 104
rect -7793 -104 -7759 -88
rect -7697 88 -7663 104
rect -7697 -104 -7663 -88
rect -7601 88 -7567 104
rect -7601 -104 -7567 -88
rect -7505 88 -7471 104
rect -7505 -104 -7471 -88
rect -7409 88 -7375 104
rect -7409 -104 -7375 -88
rect -7313 88 -7279 104
rect -7313 -104 -7279 -88
rect -7217 88 -7183 104
rect -7217 -104 -7183 -88
rect -7121 88 -7087 104
rect -7121 -104 -7087 -88
rect -7025 88 -6991 104
rect -7025 -104 -6991 -88
rect -6929 88 -6895 104
rect -6929 -104 -6895 -88
rect -6833 88 -6799 104
rect -6833 -104 -6799 -88
rect -6737 88 -6703 104
rect -6737 -104 -6703 -88
rect -6641 88 -6607 104
rect -6641 -104 -6607 -88
rect -6545 88 -6511 104
rect -6545 -104 -6511 -88
rect -6449 88 -6415 104
rect -6449 -104 -6415 -88
rect -6353 88 -6319 104
rect -6353 -104 -6319 -88
rect -6257 88 -6223 104
rect -6257 -104 -6223 -88
rect -6161 88 -6127 104
rect -6161 -104 -6127 -88
rect -6065 88 -6031 104
rect -6065 -104 -6031 -88
rect -5969 88 -5935 104
rect -5969 -104 -5935 -88
rect -5873 88 -5839 104
rect -5873 -104 -5839 -88
rect -5777 88 -5743 104
rect -5777 -104 -5743 -88
rect -5681 88 -5647 104
rect -5681 -104 -5647 -88
rect -5585 88 -5551 104
rect -5585 -104 -5551 -88
rect -5489 88 -5455 104
rect -5489 -104 -5455 -88
rect -5393 88 -5359 104
rect -5393 -104 -5359 -88
rect -5297 88 -5263 104
rect -5297 -104 -5263 -88
rect -5201 88 -5167 104
rect -5201 -104 -5167 -88
rect -5105 88 -5071 104
rect -5105 -104 -5071 -88
rect -5009 88 -4975 104
rect -5009 -104 -4975 -88
rect -4913 88 -4879 104
rect -4913 -104 -4879 -88
rect -4817 88 -4783 104
rect -4817 -104 -4783 -88
rect -4721 88 -4687 104
rect -4721 -104 -4687 -88
rect -4625 88 -4591 104
rect -4625 -104 -4591 -88
rect -4529 88 -4495 104
rect -4529 -104 -4495 -88
rect -4433 88 -4399 104
rect -4433 -104 -4399 -88
rect -4337 88 -4303 104
rect -4337 -104 -4303 -88
rect -4241 88 -4207 104
rect -4241 -104 -4207 -88
rect -4145 88 -4111 104
rect -4145 -104 -4111 -88
rect -4049 88 -4015 104
rect -4049 -104 -4015 -88
rect -3953 88 -3919 104
rect -3953 -104 -3919 -88
rect -3857 88 -3823 104
rect -3857 -104 -3823 -88
rect -3761 88 -3727 104
rect -3761 -104 -3727 -88
rect -3665 88 -3631 104
rect -3665 -104 -3631 -88
rect -3569 88 -3535 104
rect -3569 -104 -3535 -88
rect -3473 88 -3439 104
rect -3473 -104 -3439 -88
rect -3377 88 -3343 104
rect -3377 -104 -3343 -88
rect -3281 88 -3247 104
rect -3281 -104 -3247 -88
rect -3185 88 -3151 104
rect -3185 -104 -3151 -88
rect -3089 88 -3055 104
rect -3089 -104 -3055 -88
rect -2993 88 -2959 104
rect -2993 -104 -2959 -88
rect -2897 88 -2863 104
rect -2897 -104 -2863 -88
rect -2801 88 -2767 104
rect -2801 -104 -2767 -88
rect -2705 88 -2671 104
rect -2705 -104 -2671 -88
rect -2609 88 -2575 104
rect -2609 -104 -2575 -88
rect -2513 88 -2479 104
rect -2513 -104 -2479 -88
rect -2417 88 -2383 104
rect -2417 -104 -2383 -88
rect -2321 88 -2287 104
rect -2321 -104 -2287 -88
rect -2225 88 -2191 104
rect -2225 -104 -2191 -88
rect -2129 88 -2095 104
rect -2129 -104 -2095 -88
rect -2033 88 -1999 104
rect -2033 -104 -1999 -88
rect -1937 88 -1903 104
rect -1937 -104 -1903 -88
rect -1841 88 -1807 104
rect -1841 -104 -1807 -88
rect -1745 88 -1711 104
rect -1745 -104 -1711 -88
rect -1649 88 -1615 104
rect -1649 -104 -1615 -88
rect -1553 88 -1519 104
rect -1553 -104 -1519 -88
rect -1457 88 -1423 104
rect -1457 -104 -1423 -88
rect -1361 88 -1327 104
rect -1361 -104 -1327 -88
rect -1265 88 -1231 104
rect -1265 -104 -1231 -88
rect -1169 88 -1135 104
rect -1169 -104 -1135 -88
rect -1073 88 -1039 104
rect -1073 -104 -1039 -88
rect -977 88 -943 104
rect -977 -104 -943 -88
rect -881 88 -847 104
rect -881 -104 -847 -88
rect -785 88 -751 104
rect -785 -104 -751 -88
rect -689 88 -655 104
rect -689 -104 -655 -88
rect -593 88 -559 104
rect -593 -104 -559 -88
rect -497 88 -463 104
rect -497 -104 -463 -88
rect -401 88 -367 104
rect -401 -104 -367 -88
rect -305 88 -271 104
rect -305 -104 -271 -88
rect -209 88 -175 104
rect -209 -104 -175 -88
rect -113 88 -79 104
rect -113 -104 -79 -88
rect -17 88 17 104
rect -17 -104 17 -88
rect 79 88 113 104
rect 79 -104 113 -88
rect 175 88 209 104
rect 175 -104 209 -88
rect 271 88 305 104
rect 271 -104 305 -88
rect 367 88 401 104
rect 367 -104 401 -88
rect 463 88 497 104
rect 463 -104 497 -88
rect 559 88 593 104
rect 559 -104 593 -88
rect 655 88 689 104
rect 655 -104 689 -88
rect 751 88 785 104
rect 751 -104 785 -88
rect 847 88 881 104
rect 847 -104 881 -88
rect 943 88 977 104
rect 943 -104 977 -88
rect 1039 88 1073 104
rect 1039 -104 1073 -88
rect 1135 88 1169 104
rect 1135 -104 1169 -88
rect 1231 88 1265 104
rect 1231 -104 1265 -88
rect 1327 88 1361 104
rect 1327 -104 1361 -88
rect 1423 88 1457 104
rect 1423 -104 1457 -88
rect 1519 88 1553 104
rect 1519 -104 1553 -88
rect 1615 88 1649 104
rect 1615 -104 1649 -88
rect 1711 88 1745 104
rect 1711 -104 1745 -88
rect 1807 88 1841 104
rect 1807 -104 1841 -88
rect 1903 88 1937 104
rect 1903 -104 1937 -88
rect 1999 88 2033 104
rect 1999 -104 2033 -88
rect 2095 88 2129 104
rect 2095 -104 2129 -88
rect 2191 88 2225 104
rect 2191 -104 2225 -88
rect 2287 88 2321 104
rect 2287 -104 2321 -88
rect 2383 88 2417 104
rect 2383 -104 2417 -88
rect 2479 88 2513 104
rect 2479 -104 2513 -88
rect 2575 88 2609 104
rect 2575 -104 2609 -88
rect 2671 88 2705 104
rect 2671 -104 2705 -88
rect 2767 88 2801 104
rect 2767 -104 2801 -88
rect 2863 88 2897 104
rect 2863 -104 2897 -88
rect 2959 88 2993 104
rect 2959 -104 2993 -88
rect 3055 88 3089 104
rect 3055 -104 3089 -88
rect 3151 88 3185 104
rect 3151 -104 3185 -88
rect 3247 88 3281 104
rect 3247 -104 3281 -88
rect 3343 88 3377 104
rect 3343 -104 3377 -88
rect 3439 88 3473 104
rect 3439 -104 3473 -88
rect 3535 88 3569 104
rect 3535 -104 3569 -88
rect 3631 88 3665 104
rect 3631 -104 3665 -88
rect 3727 88 3761 104
rect 3727 -104 3761 -88
rect 3823 88 3857 104
rect 3823 -104 3857 -88
rect 3919 88 3953 104
rect 3919 -104 3953 -88
rect 4015 88 4049 104
rect 4015 -104 4049 -88
rect 4111 88 4145 104
rect 4111 -104 4145 -88
rect 4207 88 4241 104
rect 4207 -104 4241 -88
rect 4303 88 4337 104
rect 4303 -104 4337 -88
rect 4399 88 4433 104
rect 4399 -104 4433 -88
rect 4495 88 4529 104
rect 4495 -104 4529 -88
rect 4591 88 4625 104
rect 4591 -104 4625 -88
rect 4687 88 4721 104
rect 4687 -104 4721 -88
rect 4783 88 4817 104
rect 4783 -104 4817 -88
rect 4879 88 4913 104
rect 4879 -104 4913 -88
rect 4975 88 5009 104
rect 4975 -104 5009 -88
rect 5071 88 5105 104
rect 5071 -104 5105 -88
rect 5167 88 5201 104
rect 5167 -104 5201 -88
rect 5263 88 5297 104
rect 5263 -104 5297 -88
rect 5359 88 5393 104
rect 5359 -104 5393 -88
rect 5455 88 5489 104
rect 5455 -104 5489 -88
rect 5551 88 5585 104
rect 5551 -104 5585 -88
rect 5647 88 5681 104
rect 5647 -104 5681 -88
rect 5743 88 5777 104
rect 5743 -104 5777 -88
rect 5839 88 5873 104
rect 5839 -104 5873 -88
rect 5935 88 5969 104
rect 5935 -104 5969 -88
rect 6031 88 6065 104
rect 6031 -104 6065 -88
rect 6127 88 6161 104
rect 6127 -104 6161 -88
rect 6223 88 6257 104
rect 6223 -104 6257 -88
rect 6319 88 6353 104
rect 6319 -104 6353 -88
rect 6415 88 6449 104
rect 6415 -104 6449 -88
rect 6511 88 6545 104
rect 6511 -104 6545 -88
rect 6607 88 6641 104
rect 6607 -104 6641 -88
rect 6703 88 6737 104
rect 6703 -104 6737 -88
rect 6799 88 6833 104
rect 6799 -104 6833 -88
rect 6895 88 6929 104
rect 6895 -104 6929 -88
rect 6991 88 7025 104
rect 6991 -104 7025 -88
rect 7087 88 7121 104
rect 7087 -104 7121 -88
rect 7183 88 7217 104
rect 7183 -104 7217 -88
rect 7279 88 7313 104
rect 7279 -104 7313 -88
rect 7375 88 7409 104
rect 7375 -104 7409 -88
rect 7471 88 7505 104
rect 7471 -104 7505 -88
rect 7567 88 7601 104
rect 7567 -104 7601 -88
rect 7663 88 7697 104
rect 7663 -104 7697 -88
rect 7759 88 7793 104
rect 7759 -104 7793 -88
rect 7855 88 7889 104
rect 7855 -104 7889 -88
rect 7951 88 7985 104
rect 7951 -104 7985 -88
rect 8047 88 8081 104
rect 8047 -104 8081 -88
rect 8143 88 8177 104
rect 8143 -104 8177 -88
rect 8239 88 8273 104
rect 8239 -104 8273 -88
rect -8241 -172 -8225 -138
rect -8191 -172 -8175 -138
rect -8049 -172 -8033 -138
rect -7999 -172 -7983 -138
rect -7857 -172 -7841 -138
rect -7807 -172 -7791 -138
rect -7665 -172 -7649 -138
rect -7615 -172 -7599 -138
rect -7473 -172 -7457 -138
rect -7423 -172 -7407 -138
rect -7281 -172 -7265 -138
rect -7231 -172 -7215 -138
rect -7089 -172 -7073 -138
rect -7039 -172 -7023 -138
rect -6897 -172 -6881 -138
rect -6847 -172 -6831 -138
rect -6705 -172 -6689 -138
rect -6655 -172 -6639 -138
rect -6513 -172 -6497 -138
rect -6463 -172 -6447 -138
rect -6321 -172 -6305 -138
rect -6271 -172 -6255 -138
rect -6129 -172 -6113 -138
rect -6079 -172 -6063 -138
rect -5937 -172 -5921 -138
rect -5887 -172 -5871 -138
rect -5745 -172 -5729 -138
rect -5695 -172 -5679 -138
rect -5553 -172 -5537 -138
rect -5503 -172 -5487 -138
rect -5361 -172 -5345 -138
rect -5311 -172 -5295 -138
rect -5169 -172 -5153 -138
rect -5119 -172 -5103 -138
rect -4977 -172 -4961 -138
rect -4927 -172 -4911 -138
rect -4785 -172 -4769 -138
rect -4735 -172 -4719 -138
rect -4593 -172 -4577 -138
rect -4543 -172 -4527 -138
rect -4401 -172 -4385 -138
rect -4351 -172 -4335 -138
rect -4209 -172 -4193 -138
rect -4159 -172 -4143 -138
rect -4017 -172 -4001 -138
rect -3967 -172 -3951 -138
rect -3825 -172 -3809 -138
rect -3775 -172 -3759 -138
rect -3633 -172 -3617 -138
rect -3583 -172 -3567 -138
rect -3441 -172 -3425 -138
rect -3391 -172 -3375 -138
rect -3249 -172 -3233 -138
rect -3199 -172 -3183 -138
rect -3057 -172 -3041 -138
rect -3007 -172 -2991 -138
rect -2865 -172 -2849 -138
rect -2815 -172 -2799 -138
rect -2673 -172 -2657 -138
rect -2623 -172 -2607 -138
rect -2481 -172 -2465 -138
rect -2431 -172 -2415 -138
rect -2289 -172 -2273 -138
rect -2239 -172 -2223 -138
rect -2097 -172 -2081 -138
rect -2047 -172 -2031 -138
rect -1905 -172 -1889 -138
rect -1855 -172 -1839 -138
rect -1713 -172 -1697 -138
rect -1663 -172 -1647 -138
rect -1521 -172 -1505 -138
rect -1471 -172 -1455 -138
rect -1329 -172 -1313 -138
rect -1279 -172 -1263 -138
rect -1137 -172 -1121 -138
rect -1087 -172 -1071 -138
rect -945 -172 -929 -138
rect -895 -172 -879 -138
rect -753 -172 -737 -138
rect -703 -172 -687 -138
rect -561 -172 -545 -138
rect -511 -172 -495 -138
rect -369 -172 -353 -138
rect -319 -172 -303 -138
rect -177 -172 -161 -138
rect -127 -172 -111 -138
rect 15 -172 31 -138
rect 65 -172 81 -138
rect 207 -172 223 -138
rect 257 -172 273 -138
rect 399 -172 415 -138
rect 449 -172 465 -138
rect 591 -172 607 -138
rect 641 -172 657 -138
rect 783 -172 799 -138
rect 833 -172 849 -138
rect 975 -172 991 -138
rect 1025 -172 1041 -138
rect 1167 -172 1183 -138
rect 1217 -172 1233 -138
rect 1359 -172 1375 -138
rect 1409 -172 1425 -138
rect 1551 -172 1567 -138
rect 1601 -172 1617 -138
rect 1743 -172 1759 -138
rect 1793 -172 1809 -138
rect 1935 -172 1951 -138
rect 1985 -172 2001 -138
rect 2127 -172 2143 -138
rect 2177 -172 2193 -138
rect 2319 -172 2335 -138
rect 2369 -172 2385 -138
rect 2511 -172 2527 -138
rect 2561 -172 2577 -138
rect 2703 -172 2719 -138
rect 2753 -172 2769 -138
rect 2895 -172 2911 -138
rect 2945 -172 2961 -138
rect 3087 -172 3103 -138
rect 3137 -172 3153 -138
rect 3279 -172 3295 -138
rect 3329 -172 3345 -138
rect 3471 -172 3487 -138
rect 3521 -172 3537 -138
rect 3663 -172 3679 -138
rect 3713 -172 3729 -138
rect 3855 -172 3871 -138
rect 3905 -172 3921 -138
rect 4047 -172 4063 -138
rect 4097 -172 4113 -138
rect 4239 -172 4255 -138
rect 4289 -172 4305 -138
rect 4431 -172 4447 -138
rect 4481 -172 4497 -138
rect 4623 -172 4639 -138
rect 4673 -172 4689 -138
rect 4815 -172 4831 -138
rect 4865 -172 4881 -138
rect 5007 -172 5023 -138
rect 5057 -172 5073 -138
rect 5199 -172 5215 -138
rect 5249 -172 5265 -138
rect 5391 -172 5407 -138
rect 5441 -172 5457 -138
rect 5583 -172 5599 -138
rect 5633 -172 5649 -138
rect 5775 -172 5791 -138
rect 5825 -172 5841 -138
rect 5967 -172 5983 -138
rect 6017 -172 6033 -138
rect 6159 -172 6175 -138
rect 6209 -172 6225 -138
rect 6351 -172 6367 -138
rect 6401 -172 6417 -138
rect 6543 -172 6559 -138
rect 6593 -172 6609 -138
rect 6735 -172 6751 -138
rect 6785 -172 6801 -138
rect 6927 -172 6943 -138
rect 6977 -172 6993 -138
rect 7119 -172 7135 -138
rect 7169 -172 7185 -138
rect 7311 -172 7327 -138
rect 7361 -172 7377 -138
rect 7503 -172 7519 -138
rect 7553 -172 7569 -138
rect 7695 -172 7711 -138
rect 7745 -172 7761 -138
rect 7887 -172 7903 -138
rect 7937 -172 7953 -138
rect 8079 -172 8095 -138
rect 8129 -172 8145 -138
rect -8387 -240 -8353 -178
rect 8353 -240 8387 -178
rect -8387 -274 -8291 -240
rect 8291 -274 8387 -240
<< viali >>
rect -8129 138 -8095 172
rect -7937 138 -7903 172
rect -7745 138 -7711 172
rect -7553 138 -7519 172
rect -7361 138 -7327 172
rect -7169 138 -7135 172
rect -6977 138 -6943 172
rect -6785 138 -6751 172
rect -6593 138 -6559 172
rect -6401 138 -6367 172
rect -6209 138 -6175 172
rect -6017 138 -5983 172
rect -5825 138 -5791 172
rect -5633 138 -5599 172
rect -5441 138 -5407 172
rect -5249 138 -5215 172
rect -5057 138 -5023 172
rect -4865 138 -4831 172
rect -4673 138 -4639 172
rect -4481 138 -4447 172
rect -4289 138 -4255 172
rect -4097 138 -4063 172
rect -3905 138 -3871 172
rect -3713 138 -3679 172
rect -3521 138 -3487 172
rect -3329 138 -3295 172
rect -3137 138 -3103 172
rect -2945 138 -2911 172
rect -2753 138 -2719 172
rect -2561 138 -2527 172
rect -2369 138 -2335 172
rect -2177 138 -2143 172
rect -1985 138 -1951 172
rect -1793 138 -1759 172
rect -1601 138 -1567 172
rect -1409 138 -1375 172
rect -1217 138 -1183 172
rect -1025 138 -991 172
rect -833 138 -799 172
rect -641 138 -607 172
rect -449 138 -415 172
rect -257 138 -223 172
rect -65 138 -31 172
rect 127 138 161 172
rect 319 138 353 172
rect 511 138 545 172
rect 703 138 737 172
rect 895 138 929 172
rect 1087 138 1121 172
rect 1279 138 1313 172
rect 1471 138 1505 172
rect 1663 138 1697 172
rect 1855 138 1889 172
rect 2047 138 2081 172
rect 2239 138 2273 172
rect 2431 138 2465 172
rect 2623 138 2657 172
rect 2815 138 2849 172
rect 3007 138 3041 172
rect 3199 138 3233 172
rect 3391 138 3425 172
rect 3583 138 3617 172
rect 3775 138 3809 172
rect 3967 138 4001 172
rect 4159 138 4193 172
rect 4351 138 4385 172
rect 4543 138 4577 172
rect 4735 138 4769 172
rect 4927 138 4961 172
rect 5119 138 5153 172
rect 5311 138 5345 172
rect 5503 138 5537 172
rect 5695 138 5729 172
rect 5887 138 5921 172
rect 6079 138 6113 172
rect 6271 138 6305 172
rect 6463 138 6497 172
rect 6655 138 6689 172
rect 6847 138 6881 172
rect 7039 138 7073 172
rect 7231 138 7265 172
rect 7423 138 7457 172
rect 7615 138 7649 172
rect 7807 138 7841 172
rect 7999 138 8033 172
rect 8191 138 8225 172
rect -8273 -88 -8239 88
rect -8177 -88 -8143 88
rect -8081 -88 -8047 88
rect -7985 -88 -7951 88
rect -7889 -88 -7855 88
rect -7793 -88 -7759 88
rect -7697 -88 -7663 88
rect -7601 -88 -7567 88
rect -7505 -88 -7471 88
rect -7409 -88 -7375 88
rect -7313 -88 -7279 88
rect -7217 -88 -7183 88
rect -7121 -88 -7087 88
rect -7025 -88 -6991 88
rect -6929 -88 -6895 88
rect -6833 -88 -6799 88
rect -6737 -88 -6703 88
rect -6641 -88 -6607 88
rect -6545 -88 -6511 88
rect -6449 -88 -6415 88
rect -6353 -88 -6319 88
rect -6257 -88 -6223 88
rect -6161 -88 -6127 88
rect -6065 -88 -6031 88
rect -5969 -88 -5935 88
rect -5873 -88 -5839 88
rect -5777 -88 -5743 88
rect -5681 -88 -5647 88
rect -5585 -88 -5551 88
rect -5489 -88 -5455 88
rect -5393 -88 -5359 88
rect -5297 -88 -5263 88
rect -5201 -88 -5167 88
rect -5105 -88 -5071 88
rect -5009 -88 -4975 88
rect -4913 -88 -4879 88
rect -4817 -88 -4783 88
rect -4721 -88 -4687 88
rect -4625 -88 -4591 88
rect -4529 -88 -4495 88
rect -4433 -88 -4399 88
rect -4337 -88 -4303 88
rect -4241 -88 -4207 88
rect -4145 -88 -4111 88
rect -4049 -88 -4015 88
rect -3953 -88 -3919 88
rect -3857 -88 -3823 88
rect -3761 -88 -3727 88
rect -3665 -88 -3631 88
rect -3569 -88 -3535 88
rect -3473 -88 -3439 88
rect -3377 -88 -3343 88
rect -3281 -88 -3247 88
rect -3185 -88 -3151 88
rect -3089 -88 -3055 88
rect -2993 -88 -2959 88
rect -2897 -88 -2863 88
rect -2801 -88 -2767 88
rect -2705 -88 -2671 88
rect -2609 -88 -2575 88
rect -2513 -88 -2479 88
rect -2417 -88 -2383 88
rect -2321 -88 -2287 88
rect -2225 -88 -2191 88
rect -2129 -88 -2095 88
rect -2033 -88 -1999 88
rect -1937 -88 -1903 88
rect -1841 -88 -1807 88
rect -1745 -88 -1711 88
rect -1649 -88 -1615 88
rect -1553 -88 -1519 88
rect -1457 -88 -1423 88
rect -1361 -88 -1327 88
rect -1265 -88 -1231 88
rect -1169 -88 -1135 88
rect -1073 -88 -1039 88
rect -977 -88 -943 88
rect -881 -88 -847 88
rect -785 -88 -751 88
rect -689 -88 -655 88
rect -593 -88 -559 88
rect -497 -88 -463 88
rect -401 -88 -367 88
rect -305 -88 -271 88
rect -209 -88 -175 88
rect -113 -88 -79 88
rect -17 -88 17 88
rect 79 -88 113 88
rect 175 -88 209 88
rect 271 -88 305 88
rect 367 -88 401 88
rect 463 -88 497 88
rect 559 -88 593 88
rect 655 -88 689 88
rect 751 -88 785 88
rect 847 -88 881 88
rect 943 -88 977 88
rect 1039 -88 1073 88
rect 1135 -88 1169 88
rect 1231 -88 1265 88
rect 1327 -88 1361 88
rect 1423 -88 1457 88
rect 1519 -88 1553 88
rect 1615 -88 1649 88
rect 1711 -88 1745 88
rect 1807 -88 1841 88
rect 1903 -88 1937 88
rect 1999 -88 2033 88
rect 2095 -88 2129 88
rect 2191 -88 2225 88
rect 2287 -88 2321 88
rect 2383 -88 2417 88
rect 2479 -88 2513 88
rect 2575 -88 2609 88
rect 2671 -88 2705 88
rect 2767 -88 2801 88
rect 2863 -88 2897 88
rect 2959 -88 2993 88
rect 3055 -88 3089 88
rect 3151 -88 3185 88
rect 3247 -88 3281 88
rect 3343 -88 3377 88
rect 3439 -88 3473 88
rect 3535 -88 3569 88
rect 3631 -88 3665 88
rect 3727 -88 3761 88
rect 3823 -88 3857 88
rect 3919 -88 3953 88
rect 4015 -88 4049 88
rect 4111 -88 4145 88
rect 4207 -88 4241 88
rect 4303 -88 4337 88
rect 4399 -88 4433 88
rect 4495 -88 4529 88
rect 4591 -88 4625 88
rect 4687 -88 4721 88
rect 4783 -88 4817 88
rect 4879 -88 4913 88
rect 4975 -88 5009 88
rect 5071 -88 5105 88
rect 5167 -88 5201 88
rect 5263 -88 5297 88
rect 5359 -88 5393 88
rect 5455 -88 5489 88
rect 5551 -88 5585 88
rect 5647 -88 5681 88
rect 5743 -88 5777 88
rect 5839 -88 5873 88
rect 5935 -88 5969 88
rect 6031 -88 6065 88
rect 6127 -88 6161 88
rect 6223 -88 6257 88
rect 6319 -88 6353 88
rect 6415 -88 6449 88
rect 6511 -88 6545 88
rect 6607 -88 6641 88
rect 6703 -88 6737 88
rect 6799 -88 6833 88
rect 6895 -88 6929 88
rect 6991 -88 7025 88
rect 7087 -88 7121 88
rect 7183 -88 7217 88
rect 7279 -88 7313 88
rect 7375 -88 7409 88
rect 7471 -88 7505 88
rect 7567 -88 7601 88
rect 7663 -88 7697 88
rect 7759 -88 7793 88
rect 7855 -88 7889 88
rect 7951 -88 7985 88
rect 8047 -88 8081 88
rect 8143 -88 8177 88
rect 8239 -88 8273 88
rect -8225 -172 -8191 -138
rect -8033 -172 -7999 -138
rect -7841 -172 -7807 -138
rect -7649 -172 -7615 -138
rect -7457 -172 -7423 -138
rect -7265 -172 -7231 -138
rect -7073 -172 -7039 -138
rect -6881 -172 -6847 -138
rect -6689 -172 -6655 -138
rect -6497 -172 -6463 -138
rect -6305 -172 -6271 -138
rect -6113 -172 -6079 -138
rect -5921 -172 -5887 -138
rect -5729 -172 -5695 -138
rect -5537 -172 -5503 -138
rect -5345 -172 -5311 -138
rect -5153 -172 -5119 -138
rect -4961 -172 -4927 -138
rect -4769 -172 -4735 -138
rect -4577 -172 -4543 -138
rect -4385 -172 -4351 -138
rect -4193 -172 -4159 -138
rect -4001 -172 -3967 -138
rect -3809 -172 -3775 -138
rect -3617 -172 -3583 -138
rect -3425 -172 -3391 -138
rect -3233 -172 -3199 -138
rect -3041 -172 -3007 -138
rect -2849 -172 -2815 -138
rect -2657 -172 -2623 -138
rect -2465 -172 -2431 -138
rect -2273 -172 -2239 -138
rect -2081 -172 -2047 -138
rect -1889 -172 -1855 -138
rect -1697 -172 -1663 -138
rect -1505 -172 -1471 -138
rect -1313 -172 -1279 -138
rect -1121 -172 -1087 -138
rect -929 -172 -895 -138
rect -737 -172 -703 -138
rect -545 -172 -511 -138
rect -353 -172 -319 -138
rect -161 -172 -127 -138
rect 31 -172 65 -138
rect 223 -172 257 -138
rect 415 -172 449 -138
rect 607 -172 641 -138
rect 799 -172 833 -138
rect 991 -172 1025 -138
rect 1183 -172 1217 -138
rect 1375 -172 1409 -138
rect 1567 -172 1601 -138
rect 1759 -172 1793 -138
rect 1951 -172 1985 -138
rect 2143 -172 2177 -138
rect 2335 -172 2369 -138
rect 2527 -172 2561 -138
rect 2719 -172 2753 -138
rect 2911 -172 2945 -138
rect 3103 -172 3137 -138
rect 3295 -172 3329 -138
rect 3487 -172 3521 -138
rect 3679 -172 3713 -138
rect 3871 -172 3905 -138
rect 4063 -172 4097 -138
rect 4255 -172 4289 -138
rect 4447 -172 4481 -138
rect 4639 -172 4673 -138
rect 4831 -172 4865 -138
rect 5023 -172 5057 -138
rect 5215 -172 5249 -138
rect 5407 -172 5441 -138
rect 5599 -172 5633 -138
rect 5791 -172 5825 -138
rect 5983 -172 6017 -138
rect 6175 -172 6209 -138
rect 6367 -172 6401 -138
rect 6559 -172 6593 -138
rect 6751 -172 6785 -138
rect 6943 -172 6977 -138
rect 7135 -172 7169 -138
rect 7327 -172 7361 -138
rect 7519 -172 7553 -138
rect 7711 -172 7745 -138
rect 7903 -172 7937 -138
rect 8095 -172 8129 -138
<< metal1 >>
rect -8141 172 -8083 178
rect -8141 138 -8129 172
rect -8095 138 -8083 172
rect -8141 132 -8083 138
rect -7949 172 -7891 178
rect -7949 138 -7937 172
rect -7903 138 -7891 172
rect -7949 132 -7891 138
rect -7757 172 -7699 178
rect -7757 138 -7745 172
rect -7711 138 -7699 172
rect -7757 132 -7699 138
rect -7565 172 -7507 178
rect -7565 138 -7553 172
rect -7519 138 -7507 172
rect -7565 132 -7507 138
rect -7373 172 -7315 178
rect -7373 138 -7361 172
rect -7327 138 -7315 172
rect -7373 132 -7315 138
rect -7181 172 -7123 178
rect -7181 138 -7169 172
rect -7135 138 -7123 172
rect -7181 132 -7123 138
rect -6989 172 -6931 178
rect -6989 138 -6977 172
rect -6943 138 -6931 172
rect -6989 132 -6931 138
rect -6797 172 -6739 178
rect -6797 138 -6785 172
rect -6751 138 -6739 172
rect -6797 132 -6739 138
rect -6605 172 -6547 178
rect -6605 138 -6593 172
rect -6559 138 -6547 172
rect -6605 132 -6547 138
rect -6413 172 -6355 178
rect -6413 138 -6401 172
rect -6367 138 -6355 172
rect -6413 132 -6355 138
rect -6221 172 -6163 178
rect -6221 138 -6209 172
rect -6175 138 -6163 172
rect -6221 132 -6163 138
rect -6029 172 -5971 178
rect -6029 138 -6017 172
rect -5983 138 -5971 172
rect -6029 132 -5971 138
rect -5837 172 -5779 178
rect -5837 138 -5825 172
rect -5791 138 -5779 172
rect -5837 132 -5779 138
rect -5645 172 -5587 178
rect -5645 138 -5633 172
rect -5599 138 -5587 172
rect -5645 132 -5587 138
rect -5453 172 -5395 178
rect -5453 138 -5441 172
rect -5407 138 -5395 172
rect -5453 132 -5395 138
rect -5261 172 -5203 178
rect -5261 138 -5249 172
rect -5215 138 -5203 172
rect -5261 132 -5203 138
rect -5069 172 -5011 178
rect -5069 138 -5057 172
rect -5023 138 -5011 172
rect -5069 132 -5011 138
rect -4877 172 -4819 178
rect -4877 138 -4865 172
rect -4831 138 -4819 172
rect -4877 132 -4819 138
rect -4685 172 -4627 178
rect -4685 138 -4673 172
rect -4639 138 -4627 172
rect -4685 132 -4627 138
rect -4493 172 -4435 178
rect -4493 138 -4481 172
rect -4447 138 -4435 172
rect -4493 132 -4435 138
rect -4301 172 -4243 178
rect -4301 138 -4289 172
rect -4255 138 -4243 172
rect -4301 132 -4243 138
rect -4109 172 -4051 178
rect -4109 138 -4097 172
rect -4063 138 -4051 172
rect -4109 132 -4051 138
rect -3917 172 -3859 178
rect -3917 138 -3905 172
rect -3871 138 -3859 172
rect -3917 132 -3859 138
rect -3725 172 -3667 178
rect -3725 138 -3713 172
rect -3679 138 -3667 172
rect -3725 132 -3667 138
rect -3533 172 -3475 178
rect -3533 138 -3521 172
rect -3487 138 -3475 172
rect -3533 132 -3475 138
rect -3341 172 -3283 178
rect -3341 138 -3329 172
rect -3295 138 -3283 172
rect -3341 132 -3283 138
rect -3149 172 -3091 178
rect -3149 138 -3137 172
rect -3103 138 -3091 172
rect -3149 132 -3091 138
rect -2957 172 -2899 178
rect -2957 138 -2945 172
rect -2911 138 -2899 172
rect -2957 132 -2899 138
rect -2765 172 -2707 178
rect -2765 138 -2753 172
rect -2719 138 -2707 172
rect -2765 132 -2707 138
rect -2573 172 -2515 178
rect -2573 138 -2561 172
rect -2527 138 -2515 172
rect -2573 132 -2515 138
rect -2381 172 -2323 178
rect -2381 138 -2369 172
rect -2335 138 -2323 172
rect -2381 132 -2323 138
rect -2189 172 -2131 178
rect -2189 138 -2177 172
rect -2143 138 -2131 172
rect -2189 132 -2131 138
rect -1997 172 -1939 178
rect -1997 138 -1985 172
rect -1951 138 -1939 172
rect -1997 132 -1939 138
rect -1805 172 -1747 178
rect -1805 138 -1793 172
rect -1759 138 -1747 172
rect -1805 132 -1747 138
rect -1613 172 -1555 178
rect -1613 138 -1601 172
rect -1567 138 -1555 172
rect -1613 132 -1555 138
rect -1421 172 -1363 178
rect -1421 138 -1409 172
rect -1375 138 -1363 172
rect -1421 132 -1363 138
rect -1229 172 -1171 178
rect -1229 138 -1217 172
rect -1183 138 -1171 172
rect -1229 132 -1171 138
rect -1037 172 -979 178
rect -1037 138 -1025 172
rect -991 138 -979 172
rect -1037 132 -979 138
rect -845 172 -787 178
rect -845 138 -833 172
rect -799 138 -787 172
rect -845 132 -787 138
rect -653 172 -595 178
rect -653 138 -641 172
rect -607 138 -595 172
rect -653 132 -595 138
rect -461 172 -403 178
rect -461 138 -449 172
rect -415 138 -403 172
rect -461 132 -403 138
rect -269 172 -211 178
rect -269 138 -257 172
rect -223 138 -211 172
rect -269 132 -211 138
rect -77 172 -19 178
rect -77 138 -65 172
rect -31 138 -19 172
rect -77 132 -19 138
rect 115 172 173 178
rect 115 138 127 172
rect 161 138 173 172
rect 115 132 173 138
rect 307 172 365 178
rect 307 138 319 172
rect 353 138 365 172
rect 307 132 365 138
rect 499 172 557 178
rect 499 138 511 172
rect 545 138 557 172
rect 499 132 557 138
rect 691 172 749 178
rect 691 138 703 172
rect 737 138 749 172
rect 691 132 749 138
rect 883 172 941 178
rect 883 138 895 172
rect 929 138 941 172
rect 883 132 941 138
rect 1075 172 1133 178
rect 1075 138 1087 172
rect 1121 138 1133 172
rect 1075 132 1133 138
rect 1267 172 1325 178
rect 1267 138 1279 172
rect 1313 138 1325 172
rect 1267 132 1325 138
rect 1459 172 1517 178
rect 1459 138 1471 172
rect 1505 138 1517 172
rect 1459 132 1517 138
rect 1651 172 1709 178
rect 1651 138 1663 172
rect 1697 138 1709 172
rect 1651 132 1709 138
rect 1843 172 1901 178
rect 1843 138 1855 172
rect 1889 138 1901 172
rect 1843 132 1901 138
rect 2035 172 2093 178
rect 2035 138 2047 172
rect 2081 138 2093 172
rect 2035 132 2093 138
rect 2227 172 2285 178
rect 2227 138 2239 172
rect 2273 138 2285 172
rect 2227 132 2285 138
rect 2419 172 2477 178
rect 2419 138 2431 172
rect 2465 138 2477 172
rect 2419 132 2477 138
rect 2611 172 2669 178
rect 2611 138 2623 172
rect 2657 138 2669 172
rect 2611 132 2669 138
rect 2803 172 2861 178
rect 2803 138 2815 172
rect 2849 138 2861 172
rect 2803 132 2861 138
rect 2995 172 3053 178
rect 2995 138 3007 172
rect 3041 138 3053 172
rect 2995 132 3053 138
rect 3187 172 3245 178
rect 3187 138 3199 172
rect 3233 138 3245 172
rect 3187 132 3245 138
rect 3379 172 3437 178
rect 3379 138 3391 172
rect 3425 138 3437 172
rect 3379 132 3437 138
rect 3571 172 3629 178
rect 3571 138 3583 172
rect 3617 138 3629 172
rect 3571 132 3629 138
rect 3763 172 3821 178
rect 3763 138 3775 172
rect 3809 138 3821 172
rect 3763 132 3821 138
rect 3955 172 4013 178
rect 3955 138 3967 172
rect 4001 138 4013 172
rect 3955 132 4013 138
rect 4147 172 4205 178
rect 4147 138 4159 172
rect 4193 138 4205 172
rect 4147 132 4205 138
rect 4339 172 4397 178
rect 4339 138 4351 172
rect 4385 138 4397 172
rect 4339 132 4397 138
rect 4531 172 4589 178
rect 4531 138 4543 172
rect 4577 138 4589 172
rect 4531 132 4589 138
rect 4723 172 4781 178
rect 4723 138 4735 172
rect 4769 138 4781 172
rect 4723 132 4781 138
rect 4915 172 4973 178
rect 4915 138 4927 172
rect 4961 138 4973 172
rect 4915 132 4973 138
rect 5107 172 5165 178
rect 5107 138 5119 172
rect 5153 138 5165 172
rect 5107 132 5165 138
rect 5299 172 5357 178
rect 5299 138 5311 172
rect 5345 138 5357 172
rect 5299 132 5357 138
rect 5491 172 5549 178
rect 5491 138 5503 172
rect 5537 138 5549 172
rect 5491 132 5549 138
rect 5683 172 5741 178
rect 5683 138 5695 172
rect 5729 138 5741 172
rect 5683 132 5741 138
rect 5875 172 5933 178
rect 5875 138 5887 172
rect 5921 138 5933 172
rect 5875 132 5933 138
rect 6067 172 6125 178
rect 6067 138 6079 172
rect 6113 138 6125 172
rect 6067 132 6125 138
rect 6259 172 6317 178
rect 6259 138 6271 172
rect 6305 138 6317 172
rect 6259 132 6317 138
rect 6451 172 6509 178
rect 6451 138 6463 172
rect 6497 138 6509 172
rect 6451 132 6509 138
rect 6643 172 6701 178
rect 6643 138 6655 172
rect 6689 138 6701 172
rect 6643 132 6701 138
rect 6835 172 6893 178
rect 6835 138 6847 172
rect 6881 138 6893 172
rect 6835 132 6893 138
rect 7027 172 7085 178
rect 7027 138 7039 172
rect 7073 138 7085 172
rect 7027 132 7085 138
rect 7219 172 7277 178
rect 7219 138 7231 172
rect 7265 138 7277 172
rect 7219 132 7277 138
rect 7411 172 7469 178
rect 7411 138 7423 172
rect 7457 138 7469 172
rect 7411 132 7469 138
rect 7603 172 7661 178
rect 7603 138 7615 172
rect 7649 138 7661 172
rect 7603 132 7661 138
rect 7795 172 7853 178
rect 7795 138 7807 172
rect 7841 138 7853 172
rect 7795 132 7853 138
rect 7987 172 8045 178
rect 7987 138 7999 172
rect 8033 138 8045 172
rect 7987 132 8045 138
rect 8179 172 8237 178
rect 8179 138 8191 172
rect 8225 138 8237 172
rect 8179 132 8237 138
rect -8279 88 -8233 100
rect -8279 -88 -8273 88
rect -8239 -88 -8233 88
rect -8279 -100 -8233 -88
rect -8183 88 -8137 100
rect -8183 -88 -8177 88
rect -8143 -88 -8137 88
rect -8183 -100 -8137 -88
rect -8087 88 -8041 100
rect -8087 -88 -8081 88
rect -8047 -88 -8041 88
rect -8087 -100 -8041 -88
rect -7991 88 -7945 100
rect -7991 -88 -7985 88
rect -7951 -88 -7945 88
rect -7991 -100 -7945 -88
rect -7895 88 -7849 100
rect -7895 -88 -7889 88
rect -7855 -88 -7849 88
rect -7895 -100 -7849 -88
rect -7799 88 -7753 100
rect -7799 -88 -7793 88
rect -7759 -88 -7753 88
rect -7799 -100 -7753 -88
rect -7703 88 -7657 100
rect -7703 -88 -7697 88
rect -7663 -88 -7657 88
rect -7703 -100 -7657 -88
rect -7607 88 -7561 100
rect -7607 -88 -7601 88
rect -7567 -88 -7561 88
rect -7607 -100 -7561 -88
rect -7511 88 -7465 100
rect -7511 -88 -7505 88
rect -7471 -88 -7465 88
rect -7511 -100 -7465 -88
rect -7415 88 -7369 100
rect -7415 -88 -7409 88
rect -7375 -88 -7369 88
rect -7415 -100 -7369 -88
rect -7319 88 -7273 100
rect -7319 -88 -7313 88
rect -7279 -88 -7273 88
rect -7319 -100 -7273 -88
rect -7223 88 -7177 100
rect -7223 -88 -7217 88
rect -7183 -88 -7177 88
rect -7223 -100 -7177 -88
rect -7127 88 -7081 100
rect -7127 -88 -7121 88
rect -7087 -88 -7081 88
rect -7127 -100 -7081 -88
rect -7031 88 -6985 100
rect -7031 -88 -7025 88
rect -6991 -88 -6985 88
rect -7031 -100 -6985 -88
rect -6935 88 -6889 100
rect -6935 -88 -6929 88
rect -6895 -88 -6889 88
rect -6935 -100 -6889 -88
rect -6839 88 -6793 100
rect -6839 -88 -6833 88
rect -6799 -88 -6793 88
rect -6839 -100 -6793 -88
rect -6743 88 -6697 100
rect -6743 -88 -6737 88
rect -6703 -88 -6697 88
rect -6743 -100 -6697 -88
rect -6647 88 -6601 100
rect -6647 -88 -6641 88
rect -6607 -88 -6601 88
rect -6647 -100 -6601 -88
rect -6551 88 -6505 100
rect -6551 -88 -6545 88
rect -6511 -88 -6505 88
rect -6551 -100 -6505 -88
rect -6455 88 -6409 100
rect -6455 -88 -6449 88
rect -6415 -88 -6409 88
rect -6455 -100 -6409 -88
rect -6359 88 -6313 100
rect -6359 -88 -6353 88
rect -6319 -88 -6313 88
rect -6359 -100 -6313 -88
rect -6263 88 -6217 100
rect -6263 -88 -6257 88
rect -6223 -88 -6217 88
rect -6263 -100 -6217 -88
rect -6167 88 -6121 100
rect -6167 -88 -6161 88
rect -6127 -88 -6121 88
rect -6167 -100 -6121 -88
rect -6071 88 -6025 100
rect -6071 -88 -6065 88
rect -6031 -88 -6025 88
rect -6071 -100 -6025 -88
rect -5975 88 -5929 100
rect -5975 -88 -5969 88
rect -5935 -88 -5929 88
rect -5975 -100 -5929 -88
rect -5879 88 -5833 100
rect -5879 -88 -5873 88
rect -5839 -88 -5833 88
rect -5879 -100 -5833 -88
rect -5783 88 -5737 100
rect -5783 -88 -5777 88
rect -5743 -88 -5737 88
rect -5783 -100 -5737 -88
rect -5687 88 -5641 100
rect -5687 -88 -5681 88
rect -5647 -88 -5641 88
rect -5687 -100 -5641 -88
rect -5591 88 -5545 100
rect -5591 -88 -5585 88
rect -5551 -88 -5545 88
rect -5591 -100 -5545 -88
rect -5495 88 -5449 100
rect -5495 -88 -5489 88
rect -5455 -88 -5449 88
rect -5495 -100 -5449 -88
rect -5399 88 -5353 100
rect -5399 -88 -5393 88
rect -5359 -88 -5353 88
rect -5399 -100 -5353 -88
rect -5303 88 -5257 100
rect -5303 -88 -5297 88
rect -5263 -88 -5257 88
rect -5303 -100 -5257 -88
rect -5207 88 -5161 100
rect -5207 -88 -5201 88
rect -5167 -88 -5161 88
rect -5207 -100 -5161 -88
rect -5111 88 -5065 100
rect -5111 -88 -5105 88
rect -5071 -88 -5065 88
rect -5111 -100 -5065 -88
rect -5015 88 -4969 100
rect -5015 -88 -5009 88
rect -4975 -88 -4969 88
rect -5015 -100 -4969 -88
rect -4919 88 -4873 100
rect -4919 -88 -4913 88
rect -4879 -88 -4873 88
rect -4919 -100 -4873 -88
rect -4823 88 -4777 100
rect -4823 -88 -4817 88
rect -4783 -88 -4777 88
rect -4823 -100 -4777 -88
rect -4727 88 -4681 100
rect -4727 -88 -4721 88
rect -4687 -88 -4681 88
rect -4727 -100 -4681 -88
rect -4631 88 -4585 100
rect -4631 -88 -4625 88
rect -4591 -88 -4585 88
rect -4631 -100 -4585 -88
rect -4535 88 -4489 100
rect -4535 -88 -4529 88
rect -4495 -88 -4489 88
rect -4535 -100 -4489 -88
rect -4439 88 -4393 100
rect -4439 -88 -4433 88
rect -4399 -88 -4393 88
rect -4439 -100 -4393 -88
rect -4343 88 -4297 100
rect -4343 -88 -4337 88
rect -4303 -88 -4297 88
rect -4343 -100 -4297 -88
rect -4247 88 -4201 100
rect -4247 -88 -4241 88
rect -4207 -88 -4201 88
rect -4247 -100 -4201 -88
rect -4151 88 -4105 100
rect -4151 -88 -4145 88
rect -4111 -88 -4105 88
rect -4151 -100 -4105 -88
rect -4055 88 -4009 100
rect -4055 -88 -4049 88
rect -4015 -88 -4009 88
rect -4055 -100 -4009 -88
rect -3959 88 -3913 100
rect -3959 -88 -3953 88
rect -3919 -88 -3913 88
rect -3959 -100 -3913 -88
rect -3863 88 -3817 100
rect -3863 -88 -3857 88
rect -3823 -88 -3817 88
rect -3863 -100 -3817 -88
rect -3767 88 -3721 100
rect -3767 -88 -3761 88
rect -3727 -88 -3721 88
rect -3767 -100 -3721 -88
rect -3671 88 -3625 100
rect -3671 -88 -3665 88
rect -3631 -88 -3625 88
rect -3671 -100 -3625 -88
rect -3575 88 -3529 100
rect -3575 -88 -3569 88
rect -3535 -88 -3529 88
rect -3575 -100 -3529 -88
rect -3479 88 -3433 100
rect -3479 -88 -3473 88
rect -3439 -88 -3433 88
rect -3479 -100 -3433 -88
rect -3383 88 -3337 100
rect -3383 -88 -3377 88
rect -3343 -88 -3337 88
rect -3383 -100 -3337 -88
rect -3287 88 -3241 100
rect -3287 -88 -3281 88
rect -3247 -88 -3241 88
rect -3287 -100 -3241 -88
rect -3191 88 -3145 100
rect -3191 -88 -3185 88
rect -3151 -88 -3145 88
rect -3191 -100 -3145 -88
rect -3095 88 -3049 100
rect -3095 -88 -3089 88
rect -3055 -88 -3049 88
rect -3095 -100 -3049 -88
rect -2999 88 -2953 100
rect -2999 -88 -2993 88
rect -2959 -88 -2953 88
rect -2999 -100 -2953 -88
rect -2903 88 -2857 100
rect -2903 -88 -2897 88
rect -2863 -88 -2857 88
rect -2903 -100 -2857 -88
rect -2807 88 -2761 100
rect -2807 -88 -2801 88
rect -2767 -88 -2761 88
rect -2807 -100 -2761 -88
rect -2711 88 -2665 100
rect -2711 -88 -2705 88
rect -2671 -88 -2665 88
rect -2711 -100 -2665 -88
rect -2615 88 -2569 100
rect -2615 -88 -2609 88
rect -2575 -88 -2569 88
rect -2615 -100 -2569 -88
rect -2519 88 -2473 100
rect -2519 -88 -2513 88
rect -2479 -88 -2473 88
rect -2519 -100 -2473 -88
rect -2423 88 -2377 100
rect -2423 -88 -2417 88
rect -2383 -88 -2377 88
rect -2423 -100 -2377 -88
rect -2327 88 -2281 100
rect -2327 -88 -2321 88
rect -2287 -88 -2281 88
rect -2327 -100 -2281 -88
rect -2231 88 -2185 100
rect -2231 -88 -2225 88
rect -2191 -88 -2185 88
rect -2231 -100 -2185 -88
rect -2135 88 -2089 100
rect -2135 -88 -2129 88
rect -2095 -88 -2089 88
rect -2135 -100 -2089 -88
rect -2039 88 -1993 100
rect -2039 -88 -2033 88
rect -1999 -88 -1993 88
rect -2039 -100 -1993 -88
rect -1943 88 -1897 100
rect -1943 -88 -1937 88
rect -1903 -88 -1897 88
rect -1943 -100 -1897 -88
rect -1847 88 -1801 100
rect -1847 -88 -1841 88
rect -1807 -88 -1801 88
rect -1847 -100 -1801 -88
rect -1751 88 -1705 100
rect -1751 -88 -1745 88
rect -1711 -88 -1705 88
rect -1751 -100 -1705 -88
rect -1655 88 -1609 100
rect -1655 -88 -1649 88
rect -1615 -88 -1609 88
rect -1655 -100 -1609 -88
rect -1559 88 -1513 100
rect -1559 -88 -1553 88
rect -1519 -88 -1513 88
rect -1559 -100 -1513 -88
rect -1463 88 -1417 100
rect -1463 -88 -1457 88
rect -1423 -88 -1417 88
rect -1463 -100 -1417 -88
rect -1367 88 -1321 100
rect -1367 -88 -1361 88
rect -1327 -88 -1321 88
rect -1367 -100 -1321 -88
rect -1271 88 -1225 100
rect -1271 -88 -1265 88
rect -1231 -88 -1225 88
rect -1271 -100 -1225 -88
rect -1175 88 -1129 100
rect -1175 -88 -1169 88
rect -1135 -88 -1129 88
rect -1175 -100 -1129 -88
rect -1079 88 -1033 100
rect -1079 -88 -1073 88
rect -1039 -88 -1033 88
rect -1079 -100 -1033 -88
rect -983 88 -937 100
rect -983 -88 -977 88
rect -943 -88 -937 88
rect -983 -100 -937 -88
rect -887 88 -841 100
rect -887 -88 -881 88
rect -847 -88 -841 88
rect -887 -100 -841 -88
rect -791 88 -745 100
rect -791 -88 -785 88
rect -751 -88 -745 88
rect -791 -100 -745 -88
rect -695 88 -649 100
rect -695 -88 -689 88
rect -655 -88 -649 88
rect -695 -100 -649 -88
rect -599 88 -553 100
rect -599 -88 -593 88
rect -559 -88 -553 88
rect -599 -100 -553 -88
rect -503 88 -457 100
rect -503 -88 -497 88
rect -463 -88 -457 88
rect -503 -100 -457 -88
rect -407 88 -361 100
rect -407 -88 -401 88
rect -367 -88 -361 88
rect -407 -100 -361 -88
rect -311 88 -265 100
rect -311 -88 -305 88
rect -271 -88 -265 88
rect -311 -100 -265 -88
rect -215 88 -169 100
rect -215 -88 -209 88
rect -175 -88 -169 88
rect -215 -100 -169 -88
rect -119 88 -73 100
rect -119 -88 -113 88
rect -79 -88 -73 88
rect -119 -100 -73 -88
rect -23 88 23 100
rect -23 -88 -17 88
rect 17 -88 23 88
rect -23 -100 23 -88
rect 73 88 119 100
rect 73 -88 79 88
rect 113 -88 119 88
rect 73 -100 119 -88
rect 169 88 215 100
rect 169 -88 175 88
rect 209 -88 215 88
rect 169 -100 215 -88
rect 265 88 311 100
rect 265 -88 271 88
rect 305 -88 311 88
rect 265 -100 311 -88
rect 361 88 407 100
rect 361 -88 367 88
rect 401 -88 407 88
rect 361 -100 407 -88
rect 457 88 503 100
rect 457 -88 463 88
rect 497 -88 503 88
rect 457 -100 503 -88
rect 553 88 599 100
rect 553 -88 559 88
rect 593 -88 599 88
rect 553 -100 599 -88
rect 649 88 695 100
rect 649 -88 655 88
rect 689 -88 695 88
rect 649 -100 695 -88
rect 745 88 791 100
rect 745 -88 751 88
rect 785 -88 791 88
rect 745 -100 791 -88
rect 841 88 887 100
rect 841 -88 847 88
rect 881 -88 887 88
rect 841 -100 887 -88
rect 937 88 983 100
rect 937 -88 943 88
rect 977 -88 983 88
rect 937 -100 983 -88
rect 1033 88 1079 100
rect 1033 -88 1039 88
rect 1073 -88 1079 88
rect 1033 -100 1079 -88
rect 1129 88 1175 100
rect 1129 -88 1135 88
rect 1169 -88 1175 88
rect 1129 -100 1175 -88
rect 1225 88 1271 100
rect 1225 -88 1231 88
rect 1265 -88 1271 88
rect 1225 -100 1271 -88
rect 1321 88 1367 100
rect 1321 -88 1327 88
rect 1361 -88 1367 88
rect 1321 -100 1367 -88
rect 1417 88 1463 100
rect 1417 -88 1423 88
rect 1457 -88 1463 88
rect 1417 -100 1463 -88
rect 1513 88 1559 100
rect 1513 -88 1519 88
rect 1553 -88 1559 88
rect 1513 -100 1559 -88
rect 1609 88 1655 100
rect 1609 -88 1615 88
rect 1649 -88 1655 88
rect 1609 -100 1655 -88
rect 1705 88 1751 100
rect 1705 -88 1711 88
rect 1745 -88 1751 88
rect 1705 -100 1751 -88
rect 1801 88 1847 100
rect 1801 -88 1807 88
rect 1841 -88 1847 88
rect 1801 -100 1847 -88
rect 1897 88 1943 100
rect 1897 -88 1903 88
rect 1937 -88 1943 88
rect 1897 -100 1943 -88
rect 1993 88 2039 100
rect 1993 -88 1999 88
rect 2033 -88 2039 88
rect 1993 -100 2039 -88
rect 2089 88 2135 100
rect 2089 -88 2095 88
rect 2129 -88 2135 88
rect 2089 -100 2135 -88
rect 2185 88 2231 100
rect 2185 -88 2191 88
rect 2225 -88 2231 88
rect 2185 -100 2231 -88
rect 2281 88 2327 100
rect 2281 -88 2287 88
rect 2321 -88 2327 88
rect 2281 -100 2327 -88
rect 2377 88 2423 100
rect 2377 -88 2383 88
rect 2417 -88 2423 88
rect 2377 -100 2423 -88
rect 2473 88 2519 100
rect 2473 -88 2479 88
rect 2513 -88 2519 88
rect 2473 -100 2519 -88
rect 2569 88 2615 100
rect 2569 -88 2575 88
rect 2609 -88 2615 88
rect 2569 -100 2615 -88
rect 2665 88 2711 100
rect 2665 -88 2671 88
rect 2705 -88 2711 88
rect 2665 -100 2711 -88
rect 2761 88 2807 100
rect 2761 -88 2767 88
rect 2801 -88 2807 88
rect 2761 -100 2807 -88
rect 2857 88 2903 100
rect 2857 -88 2863 88
rect 2897 -88 2903 88
rect 2857 -100 2903 -88
rect 2953 88 2999 100
rect 2953 -88 2959 88
rect 2993 -88 2999 88
rect 2953 -100 2999 -88
rect 3049 88 3095 100
rect 3049 -88 3055 88
rect 3089 -88 3095 88
rect 3049 -100 3095 -88
rect 3145 88 3191 100
rect 3145 -88 3151 88
rect 3185 -88 3191 88
rect 3145 -100 3191 -88
rect 3241 88 3287 100
rect 3241 -88 3247 88
rect 3281 -88 3287 88
rect 3241 -100 3287 -88
rect 3337 88 3383 100
rect 3337 -88 3343 88
rect 3377 -88 3383 88
rect 3337 -100 3383 -88
rect 3433 88 3479 100
rect 3433 -88 3439 88
rect 3473 -88 3479 88
rect 3433 -100 3479 -88
rect 3529 88 3575 100
rect 3529 -88 3535 88
rect 3569 -88 3575 88
rect 3529 -100 3575 -88
rect 3625 88 3671 100
rect 3625 -88 3631 88
rect 3665 -88 3671 88
rect 3625 -100 3671 -88
rect 3721 88 3767 100
rect 3721 -88 3727 88
rect 3761 -88 3767 88
rect 3721 -100 3767 -88
rect 3817 88 3863 100
rect 3817 -88 3823 88
rect 3857 -88 3863 88
rect 3817 -100 3863 -88
rect 3913 88 3959 100
rect 3913 -88 3919 88
rect 3953 -88 3959 88
rect 3913 -100 3959 -88
rect 4009 88 4055 100
rect 4009 -88 4015 88
rect 4049 -88 4055 88
rect 4009 -100 4055 -88
rect 4105 88 4151 100
rect 4105 -88 4111 88
rect 4145 -88 4151 88
rect 4105 -100 4151 -88
rect 4201 88 4247 100
rect 4201 -88 4207 88
rect 4241 -88 4247 88
rect 4201 -100 4247 -88
rect 4297 88 4343 100
rect 4297 -88 4303 88
rect 4337 -88 4343 88
rect 4297 -100 4343 -88
rect 4393 88 4439 100
rect 4393 -88 4399 88
rect 4433 -88 4439 88
rect 4393 -100 4439 -88
rect 4489 88 4535 100
rect 4489 -88 4495 88
rect 4529 -88 4535 88
rect 4489 -100 4535 -88
rect 4585 88 4631 100
rect 4585 -88 4591 88
rect 4625 -88 4631 88
rect 4585 -100 4631 -88
rect 4681 88 4727 100
rect 4681 -88 4687 88
rect 4721 -88 4727 88
rect 4681 -100 4727 -88
rect 4777 88 4823 100
rect 4777 -88 4783 88
rect 4817 -88 4823 88
rect 4777 -100 4823 -88
rect 4873 88 4919 100
rect 4873 -88 4879 88
rect 4913 -88 4919 88
rect 4873 -100 4919 -88
rect 4969 88 5015 100
rect 4969 -88 4975 88
rect 5009 -88 5015 88
rect 4969 -100 5015 -88
rect 5065 88 5111 100
rect 5065 -88 5071 88
rect 5105 -88 5111 88
rect 5065 -100 5111 -88
rect 5161 88 5207 100
rect 5161 -88 5167 88
rect 5201 -88 5207 88
rect 5161 -100 5207 -88
rect 5257 88 5303 100
rect 5257 -88 5263 88
rect 5297 -88 5303 88
rect 5257 -100 5303 -88
rect 5353 88 5399 100
rect 5353 -88 5359 88
rect 5393 -88 5399 88
rect 5353 -100 5399 -88
rect 5449 88 5495 100
rect 5449 -88 5455 88
rect 5489 -88 5495 88
rect 5449 -100 5495 -88
rect 5545 88 5591 100
rect 5545 -88 5551 88
rect 5585 -88 5591 88
rect 5545 -100 5591 -88
rect 5641 88 5687 100
rect 5641 -88 5647 88
rect 5681 -88 5687 88
rect 5641 -100 5687 -88
rect 5737 88 5783 100
rect 5737 -88 5743 88
rect 5777 -88 5783 88
rect 5737 -100 5783 -88
rect 5833 88 5879 100
rect 5833 -88 5839 88
rect 5873 -88 5879 88
rect 5833 -100 5879 -88
rect 5929 88 5975 100
rect 5929 -88 5935 88
rect 5969 -88 5975 88
rect 5929 -100 5975 -88
rect 6025 88 6071 100
rect 6025 -88 6031 88
rect 6065 -88 6071 88
rect 6025 -100 6071 -88
rect 6121 88 6167 100
rect 6121 -88 6127 88
rect 6161 -88 6167 88
rect 6121 -100 6167 -88
rect 6217 88 6263 100
rect 6217 -88 6223 88
rect 6257 -88 6263 88
rect 6217 -100 6263 -88
rect 6313 88 6359 100
rect 6313 -88 6319 88
rect 6353 -88 6359 88
rect 6313 -100 6359 -88
rect 6409 88 6455 100
rect 6409 -88 6415 88
rect 6449 -88 6455 88
rect 6409 -100 6455 -88
rect 6505 88 6551 100
rect 6505 -88 6511 88
rect 6545 -88 6551 88
rect 6505 -100 6551 -88
rect 6601 88 6647 100
rect 6601 -88 6607 88
rect 6641 -88 6647 88
rect 6601 -100 6647 -88
rect 6697 88 6743 100
rect 6697 -88 6703 88
rect 6737 -88 6743 88
rect 6697 -100 6743 -88
rect 6793 88 6839 100
rect 6793 -88 6799 88
rect 6833 -88 6839 88
rect 6793 -100 6839 -88
rect 6889 88 6935 100
rect 6889 -88 6895 88
rect 6929 -88 6935 88
rect 6889 -100 6935 -88
rect 6985 88 7031 100
rect 6985 -88 6991 88
rect 7025 -88 7031 88
rect 6985 -100 7031 -88
rect 7081 88 7127 100
rect 7081 -88 7087 88
rect 7121 -88 7127 88
rect 7081 -100 7127 -88
rect 7177 88 7223 100
rect 7177 -88 7183 88
rect 7217 -88 7223 88
rect 7177 -100 7223 -88
rect 7273 88 7319 100
rect 7273 -88 7279 88
rect 7313 -88 7319 88
rect 7273 -100 7319 -88
rect 7369 88 7415 100
rect 7369 -88 7375 88
rect 7409 -88 7415 88
rect 7369 -100 7415 -88
rect 7465 88 7511 100
rect 7465 -88 7471 88
rect 7505 -88 7511 88
rect 7465 -100 7511 -88
rect 7561 88 7607 100
rect 7561 -88 7567 88
rect 7601 -88 7607 88
rect 7561 -100 7607 -88
rect 7657 88 7703 100
rect 7657 -88 7663 88
rect 7697 -88 7703 88
rect 7657 -100 7703 -88
rect 7753 88 7799 100
rect 7753 -88 7759 88
rect 7793 -88 7799 88
rect 7753 -100 7799 -88
rect 7849 88 7895 100
rect 7849 -88 7855 88
rect 7889 -88 7895 88
rect 7849 -100 7895 -88
rect 7945 88 7991 100
rect 7945 -88 7951 88
rect 7985 -88 7991 88
rect 7945 -100 7991 -88
rect 8041 88 8087 100
rect 8041 -88 8047 88
rect 8081 -88 8087 88
rect 8041 -100 8087 -88
rect 8137 88 8183 100
rect 8137 -88 8143 88
rect 8177 -88 8183 88
rect 8137 -100 8183 -88
rect 8233 88 8279 100
rect 8233 -88 8239 88
rect 8273 -88 8279 88
rect 8233 -100 8279 -88
rect -8237 -138 -8179 -132
rect -8237 -172 -8225 -138
rect -8191 -172 -8179 -138
rect -8237 -178 -8179 -172
rect -8045 -138 -7987 -132
rect -8045 -172 -8033 -138
rect -7999 -172 -7987 -138
rect -8045 -178 -7987 -172
rect -7853 -138 -7795 -132
rect -7853 -172 -7841 -138
rect -7807 -172 -7795 -138
rect -7853 -178 -7795 -172
rect -7661 -138 -7603 -132
rect -7661 -172 -7649 -138
rect -7615 -172 -7603 -138
rect -7661 -178 -7603 -172
rect -7469 -138 -7411 -132
rect -7469 -172 -7457 -138
rect -7423 -172 -7411 -138
rect -7469 -178 -7411 -172
rect -7277 -138 -7219 -132
rect -7277 -172 -7265 -138
rect -7231 -172 -7219 -138
rect -7277 -178 -7219 -172
rect -7085 -138 -7027 -132
rect -7085 -172 -7073 -138
rect -7039 -172 -7027 -138
rect -7085 -178 -7027 -172
rect -6893 -138 -6835 -132
rect -6893 -172 -6881 -138
rect -6847 -172 -6835 -138
rect -6893 -178 -6835 -172
rect -6701 -138 -6643 -132
rect -6701 -172 -6689 -138
rect -6655 -172 -6643 -138
rect -6701 -178 -6643 -172
rect -6509 -138 -6451 -132
rect -6509 -172 -6497 -138
rect -6463 -172 -6451 -138
rect -6509 -178 -6451 -172
rect -6317 -138 -6259 -132
rect -6317 -172 -6305 -138
rect -6271 -172 -6259 -138
rect -6317 -178 -6259 -172
rect -6125 -138 -6067 -132
rect -6125 -172 -6113 -138
rect -6079 -172 -6067 -138
rect -6125 -178 -6067 -172
rect -5933 -138 -5875 -132
rect -5933 -172 -5921 -138
rect -5887 -172 -5875 -138
rect -5933 -178 -5875 -172
rect -5741 -138 -5683 -132
rect -5741 -172 -5729 -138
rect -5695 -172 -5683 -138
rect -5741 -178 -5683 -172
rect -5549 -138 -5491 -132
rect -5549 -172 -5537 -138
rect -5503 -172 -5491 -138
rect -5549 -178 -5491 -172
rect -5357 -138 -5299 -132
rect -5357 -172 -5345 -138
rect -5311 -172 -5299 -138
rect -5357 -178 -5299 -172
rect -5165 -138 -5107 -132
rect -5165 -172 -5153 -138
rect -5119 -172 -5107 -138
rect -5165 -178 -5107 -172
rect -4973 -138 -4915 -132
rect -4973 -172 -4961 -138
rect -4927 -172 -4915 -138
rect -4973 -178 -4915 -172
rect -4781 -138 -4723 -132
rect -4781 -172 -4769 -138
rect -4735 -172 -4723 -138
rect -4781 -178 -4723 -172
rect -4589 -138 -4531 -132
rect -4589 -172 -4577 -138
rect -4543 -172 -4531 -138
rect -4589 -178 -4531 -172
rect -4397 -138 -4339 -132
rect -4397 -172 -4385 -138
rect -4351 -172 -4339 -138
rect -4397 -178 -4339 -172
rect -4205 -138 -4147 -132
rect -4205 -172 -4193 -138
rect -4159 -172 -4147 -138
rect -4205 -178 -4147 -172
rect -4013 -138 -3955 -132
rect -4013 -172 -4001 -138
rect -3967 -172 -3955 -138
rect -4013 -178 -3955 -172
rect -3821 -138 -3763 -132
rect -3821 -172 -3809 -138
rect -3775 -172 -3763 -138
rect -3821 -178 -3763 -172
rect -3629 -138 -3571 -132
rect -3629 -172 -3617 -138
rect -3583 -172 -3571 -138
rect -3629 -178 -3571 -172
rect -3437 -138 -3379 -132
rect -3437 -172 -3425 -138
rect -3391 -172 -3379 -138
rect -3437 -178 -3379 -172
rect -3245 -138 -3187 -132
rect -3245 -172 -3233 -138
rect -3199 -172 -3187 -138
rect -3245 -178 -3187 -172
rect -3053 -138 -2995 -132
rect -3053 -172 -3041 -138
rect -3007 -172 -2995 -138
rect -3053 -178 -2995 -172
rect -2861 -138 -2803 -132
rect -2861 -172 -2849 -138
rect -2815 -172 -2803 -138
rect -2861 -178 -2803 -172
rect -2669 -138 -2611 -132
rect -2669 -172 -2657 -138
rect -2623 -172 -2611 -138
rect -2669 -178 -2611 -172
rect -2477 -138 -2419 -132
rect -2477 -172 -2465 -138
rect -2431 -172 -2419 -138
rect -2477 -178 -2419 -172
rect -2285 -138 -2227 -132
rect -2285 -172 -2273 -138
rect -2239 -172 -2227 -138
rect -2285 -178 -2227 -172
rect -2093 -138 -2035 -132
rect -2093 -172 -2081 -138
rect -2047 -172 -2035 -138
rect -2093 -178 -2035 -172
rect -1901 -138 -1843 -132
rect -1901 -172 -1889 -138
rect -1855 -172 -1843 -138
rect -1901 -178 -1843 -172
rect -1709 -138 -1651 -132
rect -1709 -172 -1697 -138
rect -1663 -172 -1651 -138
rect -1709 -178 -1651 -172
rect -1517 -138 -1459 -132
rect -1517 -172 -1505 -138
rect -1471 -172 -1459 -138
rect -1517 -178 -1459 -172
rect -1325 -138 -1267 -132
rect -1325 -172 -1313 -138
rect -1279 -172 -1267 -138
rect -1325 -178 -1267 -172
rect -1133 -138 -1075 -132
rect -1133 -172 -1121 -138
rect -1087 -172 -1075 -138
rect -1133 -178 -1075 -172
rect -941 -138 -883 -132
rect -941 -172 -929 -138
rect -895 -172 -883 -138
rect -941 -178 -883 -172
rect -749 -138 -691 -132
rect -749 -172 -737 -138
rect -703 -172 -691 -138
rect -749 -178 -691 -172
rect -557 -138 -499 -132
rect -557 -172 -545 -138
rect -511 -172 -499 -138
rect -557 -178 -499 -172
rect -365 -138 -307 -132
rect -365 -172 -353 -138
rect -319 -172 -307 -138
rect -365 -178 -307 -172
rect -173 -138 -115 -132
rect -173 -172 -161 -138
rect -127 -172 -115 -138
rect -173 -178 -115 -172
rect 19 -138 77 -132
rect 19 -172 31 -138
rect 65 -172 77 -138
rect 19 -178 77 -172
rect 211 -138 269 -132
rect 211 -172 223 -138
rect 257 -172 269 -138
rect 211 -178 269 -172
rect 403 -138 461 -132
rect 403 -172 415 -138
rect 449 -172 461 -138
rect 403 -178 461 -172
rect 595 -138 653 -132
rect 595 -172 607 -138
rect 641 -172 653 -138
rect 595 -178 653 -172
rect 787 -138 845 -132
rect 787 -172 799 -138
rect 833 -172 845 -138
rect 787 -178 845 -172
rect 979 -138 1037 -132
rect 979 -172 991 -138
rect 1025 -172 1037 -138
rect 979 -178 1037 -172
rect 1171 -138 1229 -132
rect 1171 -172 1183 -138
rect 1217 -172 1229 -138
rect 1171 -178 1229 -172
rect 1363 -138 1421 -132
rect 1363 -172 1375 -138
rect 1409 -172 1421 -138
rect 1363 -178 1421 -172
rect 1555 -138 1613 -132
rect 1555 -172 1567 -138
rect 1601 -172 1613 -138
rect 1555 -178 1613 -172
rect 1747 -138 1805 -132
rect 1747 -172 1759 -138
rect 1793 -172 1805 -138
rect 1747 -178 1805 -172
rect 1939 -138 1997 -132
rect 1939 -172 1951 -138
rect 1985 -172 1997 -138
rect 1939 -178 1997 -172
rect 2131 -138 2189 -132
rect 2131 -172 2143 -138
rect 2177 -172 2189 -138
rect 2131 -178 2189 -172
rect 2323 -138 2381 -132
rect 2323 -172 2335 -138
rect 2369 -172 2381 -138
rect 2323 -178 2381 -172
rect 2515 -138 2573 -132
rect 2515 -172 2527 -138
rect 2561 -172 2573 -138
rect 2515 -178 2573 -172
rect 2707 -138 2765 -132
rect 2707 -172 2719 -138
rect 2753 -172 2765 -138
rect 2707 -178 2765 -172
rect 2899 -138 2957 -132
rect 2899 -172 2911 -138
rect 2945 -172 2957 -138
rect 2899 -178 2957 -172
rect 3091 -138 3149 -132
rect 3091 -172 3103 -138
rect 3137 -172 3149 -138
rect 3091 -178 3149 -172
rect 3283 -138 3341 -132
rect 3283 -172 3295 -138
rect 3329 -172 3341 -138
rect 3283 -178 3341 -172
rect 3475 -138 3533 -132
rect 3475 -172 3487 -138
rect 3521 -172 3533 -138
rect 3475 -178 3533 -172
rect 3667 -138 3725 -132
rect 3667 -172 3679 -138
rect 3713 -172 3725 -138
rect 3667 -178 3725 -172
rect 3859 -138 3917 -132
rect 3859 -172 3871 -138
rect 3905 -172 3917 -138
rect 3859 -178 3917 -172
rect 4051 -138 4109 -132
rect 4051 -172 4063 -138
rect 4097 -172 4109 -138
rect 4051 -178 4109 -172
rect 4243 -138 4301 -132
rect 4243 -172 4255 -138
rect 4289 -172 4301 -138
rect 4243 -178 4301 -172
rect 4435 -138 4493 -132
rect 4435 -172 4447 -138
rect 4481 -172 4493 -138
rect 4435 -178 4493 -172
rect 4627 -138 4685 -132
rect 4627 -172 4639 -138
rect 4673 -172 4685 -138
rect 4627 -178 4685 -172
rect 4819 -138 4877 -132
rect 4819 -172 4831 -138
rect 4865 -172 4877 -138
rect 4819 -178 4877 -172
rect 5011 -138 5069 -132
rect 5011 -172 5023 -138
rect 5057 -172 5069 -138
rect 5011 -178 5069 -172
rect 5203 -138 5261 -132
rect 5203 -172 5215 -138
rect 5249 -172 5261 -138
rect 5203 -178 5261 -172
rect 5395 -138 5453 -132
rect 5395 -172 5407 -138
rect 5441 -172 5453 -138
rect 5395 -178 5453 -172
rect 5587 -138 5645 -132
rect 5587 -172 5599 -138
rect 5633 -172 5645 -138
rect 5587 -178 5645 -172
rect 5779 -138 5837 -132
rect 5779 -172 5791 -138
rect 5825 -172 5837 -138
rect 5779 -178 5837 -172
rect 5971 -138 6029 -132
rect 5971 -172 5983 -138
rect 6017 -172 6029 -138
rect 5971 -178 6029 -172
rect 6163 -138 6221 -132
rect 6163 -172 6175 -138
rect 6209 -172 6221 -138
rect 6163 -178 6221 -172
rect 6355 -138 6413 -132
rect 6355 -172 6367 -138
rect 6401 -172 6413 -138
rect 6355 -178 6413 -172
rect 6547 -138 6605 -132
rect 6547 -172 6559 -138
rect 6593 -172 6605 -138
rect 6547 -178 6605 -172
rect 6739 -138 6797 -132
rect 6739 -172 6751 -138
rect 6785 -172 6797 -138
rect 6739 -178 6797 -172
rect 6931 -138 6989 -132
rect 6931 -172 6943 -138
rect 6977 -172 6989 -138
rect 6931 -178 6989 -172
rect 7123 -138 7181 -132
rect 7123 -172 7135 -138
rect 7169 -172 7181 -138
rect 7123 -178 7181 -172
rect 7315 -138 7373 -132
rect 7315 -172 7327 -138
rect 7361 -172 7373 -138
rect 7315 -178 7373 -172
rect 7507 -138 7565 -132
rect 7507 -172 7519 -138
rect 7553 -172 7565 -138
rect 7507 -178 7565 -172
rect 7699 -138 7757 -132
rect 7699 -172 7711 -138
rect 7745 -172 7757 -138
rect 7699 -178 7757 -172
rect 7891 -138 7949 -132
rect 7891 -172 7903 -138
rect 7937 -172 7949 -138
rect 7891 -178 7949 -172
rect 8083 -138 8141 -132
rect 8083 -172 8095 -138
rect 8129 -172 8141 -138
rect 8083 -178 8141 -172
<< properties >>
string FIXED_BBOX -8370 -257 8370 257
string gencell sky130_fd_pr__nfet_01v8_lvt
string library sky130
string parameters w 1.0 l 0.15 m 1 nf 172 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
