magic
tech sky130A
magscale 1 2
timestamp 1662478139
<< metal3 >>
rect -2650 10522 2649 10550
rect -2650 5378 2565 10522
rect 2629 5378 2649 10522
rect -2650 5350 2649 5378
rect -2650 5222 2649 5250
rect -2650 78 2565 5222
rect 2629 78 2649 5222
rect -2650 50 2649 78
rect -2650 -78 2649 -50
rect -2650 -5222 2565 -78
rect 2629 -5222 2649 -78
rect -2650 -5250 2649 -5222
rect -2650 -5378 2649 -5350
rect -2650 -10522 2565 -5378
rect 2629 -10522 2649 -5378
rect -2650 -10550 2649 -10522
<< via3 >>
rect 2565 5378 2629 10522
rect 2565 78 2629 5222
rect 2565 -5222 2629 -78
rect 2565 -10522 2629 -5378
<< mimcap >>
rect -2550 10410 2450 10450
rect -2550 5490 -2510 10410
rect 2410 5490 2450 10410
rect -2550 5450 2450 5490
rect -2550 5110 2450 5150
rect -2550 190 -2510 5110
rect 2410 190 2450 5110
rect -2550 150 2450 190
rect -2550 -190 2450 -150
rect -2550 -5110 -2510 -190
rect 2410 -5110 2450 -190
rect -2550 -5150 2450 -5110
rect -2550 -5490 2450 -5450
rect -2550 -10410 -2510 -5490
rect 2410 -10410 2450 -5490
rect -2550 -10450 2450 -10410
<< mimcapcontact >>
rect -2510 5490 2410 10410
rect -2510 190 2410 5110
rect -2510 -5110 2410 -190
rect -2510 -10410 2410 -5490
<< metal4 >>
rect -102 10411 2 10600
rect 2518 10538 2622 10600
rect 2518 10522 2645 10538
rect -2511 10410 2411 10411
rect -2511 5490 -2510 10410
rect 2410 5490 2411 10410
rect -2511 5489 2411 5490
rect -102 5111 2 5489
rect 2518 5378 2565 10522
rect 2629 5378 2645 10522
rect 2518 5362 2645 5378
rect 2518 5238 2622 5362
rect 2518 5222 2645 5238
rect -2511 5110 2411 5111
rect -2511 190 -2510 5110
rect 2410 190 2411 5110
rect -2511 189 2411 190
rect -102 -189 2 189
rect 2518 78 2565 5222
rect 2629 78 2645 5222
rect 2518 62 2645 78
rect 2518 -62 2622 62
rect 2518 -78 2645 -62
rect -2511 -190 2411 -189
rect -2511 -5110 -2510 -190
rect 2410 -5110 2411 -190
rect -2511 -5111 2411 -5110
rect -102 -5489 2 -5111
rect 2518 -5222 2565 -78
rect 2629 -5222 2645 -78
rect 2518 -5238 2645 -5222
rect 2518 -5362 2622 -5238
rect 2518 -5378 2645 -5362
rect -2511 -5490 2411 -5489
rect -2511 -10410 -2510 -5490
rect 2410 -10410 2411 -5490
rect -2511 -10411 2411 -10410
rect -102 -10600 2 -10411
rect 2518 -10522 2565 -5378
rect 2629 -10522 2645 -5378
rect 2518 -10538 2645 -10522
rect 2518 -10600 2622 -10538
<< properties >>
string FIXED_BBOX -2650 5350 2550 10550
string gencell sky130_fd_pr__cap_mim_m3_1
string library sky130
string parameters w 25.0 l 25.0 val 1.269k carea 2.00 cperi 0.19 nx 1 ny 4 dummy 0 square 0 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 1 tconnect 1 ccov 100
<< end >>
