magic
tech sky130A
magscale 1 2
timestamp 1661639644
<< nwell >>
rect -1273 -2973 1273 2973
<< pmoslvt >>
rect -1077 1554 -977 2754
rect -919 1554 -819 2754
rect -761 1554 -661 2754
rect -603 1554 -503 2754
rect -445 1554 -345 2754
rect -287 1554 -187 2754
rect -129 1554 -29 2754
rect 29 1554 129 2754
rect 187 1554 287 2754
rect 345 1554 445 2754
rect 503 1554 603 2754
rect 661 1554 761 2754
rect 819 1554 919 2754
rect 977 1554 1077 2754
rect -1077 118 -977 1318
rect -919 118 -819 1318
rect -761 118 -661 1318
rect -603 118 -503 1318
rect -445 118 -345 1318
rect -287 118 -187 1318
rect -129 118 -29 1318
rect 29 118 129 1318
rect 187 118 287 1318
rect 345 118 445 1318
rect 503 118 603 1318
rect 661 118 761 1318
rect 819 118 919 1318
rect 977 118 1077 1318
rect -1077 -1318 -977 -118
rect -919 -1318 -819 -118
rect -761 -1318 -661 -118
rect -603 -1318 -503 -118
rect -445 -1318 -345 -118
rect -287 -1318 -187 -118
rect -129 -1318 -29 -118
rect 29 -1318 129 -118
rect 187 -1318 287 -118
rect 345 -1318 445 -118
rect 503 -1318 603 -118
rect 661 -1318 761 -118
rect 819 -1318 919 -118
rect 977 -1318 1077 -118
rect -1077 -2754 -977 -1554
rect -919 -2754 -819 -1554
rect -761 -2754 -661 -1554
rect -603 -2754 -503 -1554
rect -445 -2754 -345 -1554
rect -287 -2754 -187 -1554
rect -129 -2754 -29 -1554
rect 29 -2754 129 -1554
rect 187 -2754 287 -1554
rect 345 -2754 445 -1554
rect 503 -2754 603 -1554
rect 661 -2754 761 -1554
rect 819 -2754 919 -1554
rect 977 -2754 1077 -1554
<< pdiff >>
rect -1135 2742 -1077 2754
rect -1135 1566 -1123 2742
rect -1089 1566 -1077 2742
rect -1135 1554 -1077 1566
rect -977 2742 -919 2754
rect -977 1566 -965 2742
rect -931 1566 -919 2742
rect -977 1554 -919 1566
rect -819 2742 -761 2754
rect -819 1566 -807 2742
rect -773 1566 -761 2742
rect -819 1554 -761 1566
rect -661 2742 -603 2754
rect -661 1566 -649 2742
rect -615 1566 -603 2742
rect -661 1554 -603 1566
rect -503 2742 -445 2754
rect -503 1566 -491 2742
rect -457 1566 -445 2742
rect -503 1554 -445 1566
rect -345 2742 -287 2754
rect -345 1566 -333 2742
rect -299 1566 -287 2742
rect -345 1554 -287 1566
rect -187 2742 -129 2754
rect -187 1566 -175 2742
rect -141 1566 -129 2742
rect -187 1554 -129 1566
rect -29 2742 29 2754
rect -29 1566 -17 2742
rect 17 1566 29 2742
rect -29 1554 29 1566
rect 129 2742 187 2754
rect 129 1566 141 2742
rect 175 1566 187 2742
rect 129 1554 187 1566
rect 287 2742 345 2754
rect 287 1566 299 2742
rect 333 1566 345 2742
rect 287 1554 345 1566
rect 445 2742 503 2754
rect 445 1566 457 2742
rect 491 1566 503 2742
rect 445 1554 503 1566
rect 603 2742 661 2754
rect 603 1566 615 2742
rect 649 1566 661 2742
rect 603 1554 661 1566
rect 761 2742 819 2754
rect 761 1566 773 2742
rect 807 1566 819 2742
rect 761 1554 819 1566
rect 919 2742 977 2754
rect 919 1566 931 2742
rect 965 1566 977 2742
rect 919 1554 977 1566
rect 1077 2742 1135 2754
rect 1077 1566 1089 2742
rect 1123 1566 1135 2742
rect 1077 1554 1135 1566
rect -1135 1306 -1077 1318
rect -1135 130 -1123 1306
rect -1089 130 -1077 1306
rect -1135 118 -1077 130
rect -977 1306 -919 1318
rect -977 130 -965 1306
rect -931 130 -919 1306
rect -977 118 -919 130
rect -819 1306 -761 1318
rect -819 130 -807 1306
rect -773 130 -761 1306
rect -819 118 -761 130
rect -661 1306 -603 1318
rect -661 130 -649 1306
rect -615 130 -603 1306
rect -661 118 -603 130
rect -503 1306 -445 1318
rect -503 130 -491 1306
rect -457 130 -445 1306
rect -503 118 -445 130
rect -345 1306 -287 1318
rect -345 130 -333 1306
rect -299 130 -287 1306
rect -345 118 -287 130
rect -187 1306 -129 1318
rect -187 130 -175 1306
rect -141 130 -129 1306
rect -187 118 -129 130
rect -29 1306 29 1318
rect -29 130 -17 1306
rect 17 130 29 1306
rect -29 118 29 130
rect 129 1306 187 1318
rect 129 130 141 1306
rect 175 130 187 1306
rect 129 118 187 130
rect 287 1306 345 1318
rect 287 130 299 1306
rect 333 130 345 1306
rect 287 118 345 130
rect 445 1306 503 1318
rect 445 130 457 1306
rect 491 130 503 1306
rect 445 118 503 130
rect 603 1306 661 1318
rect 603 130 615 1306
rect 649 130 661 1306
rect 603 118 661 130
rect 761 1306 819 1318
rect 761 130 773 1306
rect 807 130 819 1306
rect 761 118 819 130
rect 919 1306 977 1318
rect 919 130 931 1306
rect 965 130 977 1306
rect 919 118 977 130
rect 1077 1306 1135 1318
rect 1077 130 1089 1306
rect 1123 130 1135 1306
rect 1077 118 1135 130
rect -1135 -130 -1077 -118
rect -1135 -1306 -1123 -130
rect -1089 -1306 -1077 -130
rect -1135 -1318 -1077 -1306
rect -977 -130 -919 -118
rect -977 -1306 -965 -130
rect -931 -1306 -919 -130
rect -977 -1318 -919 -1306
rect -819 -130 -761 -118
rect -819 -1306 -807 -130
rect -773 -1306 -761 -130
rect -819 -1318 -761 -1306
rect -661 -130 -603 -118
rect -661 -1306 -649 -130
rect -615 -1306 -603 -130
rect -661 -1318 -603 -1306
rect -503 -130 -445 -118
rect -503 -1306 -491 -130
rect -457 -1306 -445 -130
rect -503 -1318 -445 -1306
rect -345 -130 -287 -118
rect -345 -1306 -333 -130
rect -299 -1306 -287 -130
rect -345 -1318 -287 -1306
rect -187 -130 -129 -118
rect -187 -1306 -175 -130
rect -141 -1306 -129 -130
rect -187 -1318 -129 -1306
rect -29 -130 29 -118
rect -29 -1306 -17 -130
rect 17 -1306 29 -130
rect -29 -1318 29 -1306
rect 129 -130 187 -118
rect 129 -1306 141 -130
rect 175 -1306 187 -130
rect 129 -1318 187 -1306
rect 287 -130 345 -118
rect 287 -1306 299 -130
rect 333 -1306 345 -130
rect 287 -1318 345 -1306
rect 445 -130 503 -118
rect 445 -1306 457 -130
rect 491 -1306 503 -130
rect 445 -1318 503 -1306
rect 603 -130 661 -118
rect 603 -1306 615 -130
rect 649 -1306 661 -130
rect 603 -1318 661 -1306
rect 761 -130 819 -118
rect 761 -1306 773 -130
rect 807 -1306 819 -130
rect 761 -1318 819 -1306
rect 919 -130 977 -118
rect 919 -1306 931 -130
rect 965 -1306 977 -130
rect 919 -1318 977 -1306
rect 1077 -130 1135 -118
rect 1077 -1306 1089 -130
rect 1123 -1306 1135 -130
rect 1077 -1318 1135 -1306
rect -1135 -1566 -1077 -1554
rect -1135 -2742 -1123 -1566
rect -1089 -2742 -1077 -1566
rect -1135 -2754 -1077 -2742
rect -977 -1566 -919 -1554
rect -977 -2742 -965 -1566
rect -931 -2742 -919 -1566
rect -977 -2754 -919 -2742
rect -819 -1566 -761 -1554
rect -819 -2742 -807 -1566
rect -773 -2742 -761 -1566
rect -819 -2754 -761 -2742
rect -661 -1566 -603 -1554
rect -661 -2742 -649 -1566
rect -615 -2742 -603 -1566
rect -661 -2754 -603 -2742
rect -503 -1566 -445 -1554
rect -503 -2742 -491 -1566
rect -457 -2742 -445 -1566
rect -503 -2754 -445 -2742
rect -345 -1566 -287 -1554
rect -345 -2742 -333 -1566
rect -299 -2742 -287 -1566
rect -345 -2754 -287 -2742
rect -187 -1566 -129 -1554
rect -187 -2742 -175 -1566
rect -141 -2742 -129 -1566
rect -187 -2754 -129 -2742
rect -29 -1566 29 -1554
rect -29 -2742 -17 -1566
rect 17 -2742 29 -1566
rect -29 -2754 29 -2742
rect 129 -1566 187 -1554
rect 129 -2742 141 -1566
rect 175 -2742 187 -1566
rect 129 -2754 187 -2742
rect 287 -1566 345 -1554
rect 287 -2742 299 -1566
rect 333 -2742 345 -1566
rect 287 -2754 345 -2742
rect 445 -1566 503 -1554
rect 445 -2742 457 -1566
rect 491 -2742 503 -1566
rect 445 -2754 503 -2742
rect 603 -1566 661 -1554
rect 603 -2742 615 -1566
rect 649 -2742 661 -1566
rect 603 -2754 661 -2742
rect 761 -1566 819 -1554
rect 761 -2742 773 -1566
rect 807 -2742 819 -1566
rect 761 -2754 819 -2742
rect 919 -1566 977 -1554
rect 919 -2742 931 -1566
rect 965 -2742 977 -1566
rect 919 -2754 977 -2742
rect 1077 -1566 1135 -1554
rect 1077 -2742 1089 -1566
rect 1123 -2742 1135 -1566
rect 1077 -2754 1135 -2742
<< pdiffc >>
rect -1123 1566 -1089 2742
rect -965 1566 -931 2742
rect -807 1566 -773 2742
rect -649 1566 -615 2742
rect -491 1566 -457 2742
rect -333 1566 -299 2742
rect -175 1566 -141 2742
rect -17 1566 17 2742
rect 141 1566 175 2742
rect 299 1566 333 2742
rect 457 1566 491 2742
rect 615 1566 649 2742
rect 773 1566 807 2742
rect 931 1566 965 2742
rect 1089 1566 1123 2742
rect -1123 130 -1089 1306
rect -965 130 -931 1306
rect -807 130 -773 1306
rect -649 130 -615 1306
rect -491 130 -457 1306
rect -333 130 -299 1306
rect -175 130 -141 1306
rect -17 130 17 1306
rect 141 130 175 1306
rect 299 130 333 1306
rect 457 130 491 1306
rect 615 130 649 1306
rect 773 130 807 1306
rect 931 130 965 1306
rect 1089 130 1123 1306
rect -1123 -1306 -1089 -130
rect -965 -1306 -931 -130
rect -807 -1306 -773 -130
rect -649 -1306 -615 -130
rect -491 -1306 -457 -130
rect -333 -1306 -299 -130
rect -175 -1306 -141 -130
rect -17 -1306 17 -130
rect 141 -1306 175 -130
rect 299 -1306 333 -130
rect 457 -1306 491 -130
rect 615 -1306 649 -130
rect 773 -1306 807 -130
rect 931 -1306 965 -130
rect 1089 -1306 1123 -130
rect -1123 -2742 -1089 -1566
rect -965 -2742 -931 -1566
rect -807 -2742 -773 -1566
rect -649 -2742 -615 -1566
rect -491 -2742 -457 -1566
rect -333 -2742 -299 -1566
rect -175 -2742 -141 -1566
rect -17 -2742 17 -1566
rect 141 -2742 175 -1566
rect 299 -2742 333 -1566
rect 457 -2742 491 -1566
rect 615 -2742 649 -1566
rect 773 -2742 807 -1566
rect 931 -2742 965 -1566
rect 1089 -2742 1123 -1566
<< nsubdiff >>
rect -1237 2903 -1141 2937
rect 1141 2903 1237 2937
rect -1237 2841 -1203 2903
rect 1203 2841 1237 2903
rect -1237 -2903 -1203 -2841
rect 1203 -2903 1237 -2841
rect -1237 -2937 -1141 -2903
rect 1141 -2937 1237 -2903
<< nsubdiffcont >>
rect -1141 2903 1141 2937
rect -1237 -2841 -1203 2841
rect 1203 -2841 1237 2841
rect -1141 -2937 1141 -2903
<< poly >>
rect -1077 2835 -977 2851
rect -1077 2801 -1061 2835
rect -993 2801 -977 2835
rect -1077 2754 -977 2801
rect -919 2835 -819 2851
rect -919 2801 -903 2835
rect -835 2801 -819 2835
rect -919 2754 -819 2801
rect -761 2835 -661 2851
rect -761 2801 -745 2835
rect -677 2801 -661 2835
rect -761 2754 -661 2801
rect -603 2835 -503 2851
rect -603 2801 -587 2835
rect -519 2801 -503 2835
rect -603 2754 -503 2801
rect -445 2835 -345 2851
rect -445 2801 -429 2835
rect -361 2801 -345 2835
rect -445 2754 -345 2801
rect -287 2835 -187 2851
rect -287 2801 -271 2835
rect -203 2801 -187 2835
rect -287 2754 -187 2801
rect -129 2835 -29 2851
rect -129 2801 -113 2835
rect -45 2801 -29 2835
rect -129 2754 -29 2801
rect 29 2835 129 2851
rect 29 2801 45 2835
rect 113 2801 129 2835
rect 29 2754 129 2801
rect 187 2835 287 2851
rect 187 2801 203 2835
rect 271 2801 287 2835
rect 187 2754 287 2801
rect 345 2835 445 2851
rect 345 2801 361 2835
rect 429 2801 445 2835
rect 345 2754 445 2801
rect 503 2835 603 2851
rect 503 2801 519 2835
rect 587 2801 603 2835
rect 503 2754 603 2801
rect 661 2835 761 2851
rect 661 2801 677 2835
rect 745 2801 761 2835
rect 661 2754 761 2801
rect 819 2835 919 2851
rect 819 2801 835 2835
rect 903 2801 919 2835
rect 819 2754 919 2801
rect 977 2835 1077 2851
rect 977 2801 993 2835
rect 1061 2801 1077 2835
rect 977 2754 1077 2801
rect -1077 1507 -977 1554
rect -1077 1473 -1061 1507
rect -993 1473 -977 1507
rect -1077 1457 -977 1473
rect -919 1507 -819 1554
rect -919 1473 -903 1507
rect -835 1473 -819 1507
rect -919 1457 -819 1473
rect -761 1507 -661 1554
rect -761 1473 -745 1507
rect -677 1473 -661 1507
rect -761 1457 -661 1473
rect -603 1507 -503 1554
rect -603 1473 -587 1507
rect -519 1473 -503 1507
rect -603 1457 -503 1473
rect -445 1507 -345 1554
rect -445 1473 -429 1507
rect -361 1473 -345 1507
rect -445 1457 -345 1473
rect -287 1507 -187 1554
rect -287 1473 -271 1507
rect -203 1473 -187 1507
rect -287 1457 -187 1473
rect -129 1507 -29 1554
rect -129 1473 -113 1507
rect -45 1473 -29 1507
rect -129 1457 -29 1473
rect 29 1507 129 1554
rect 29 1473 45 1507
rect 113 1473 129 1507
rect 29 1457 129 1473
rect 187 1507 287 1554
rect 187 1473 203 1507
rect 271 1473 287 1507
rect 187 1457 287 1473
rect 345 1507 445 1554
rect 345 1473 361 1507
rect 429 1473 445 1507
rect 345 1457 445 1473
rect 503 1507 603 1554
rect 503 1473 519 1507
rect 587 1473 603 1507
rect 503 1457 603 1473
rect 661 1507 761 1554
rect 661 1473 677 1507
rect 745 1473 761 1507
rect 661 1457 761 1473
rect 819 1507 919 1554
rect 819 1473 835 1507
rect 903 1473 919 1507
rect 819 1457 919 1473
rect 977 1507 1077 1554
rect 977 1473 993 1507
rect 1061 1473 1077 1507
rect 977 1457 1077 1473
rect -1077 1399 -977 1415
rect -1077 1365 -1061 1399
rect -993 1365 -977 1399
rect -1077 1318 -977 1365
rect -919 1399 -819 1415
rect -919 1365 -903 1399
rect -835 1365 -819 1399
rect -919 1318 -819 1365
rect -761 1399 -661 1415
rect -761 1365 -745 1399
rect -677 1365 -661 1399
rect -761 1318 -661 1365
rect -603 1399 -503 1415
rect -603 1365 -587 1399
rect -519 1365 -503 1399
rect -603 1318 -503 1365
rect -445 1399 -345 1415
rect -445 1365 -429 1399
rect -361 1365 -345 1399
rect -445 1318 -345 1365
rect -287 1399 -187 1415
rect -287 1365 -271 1399
rect -203 1365 -187 1399
rect -287 1318 -187 1365
rect -129 1399 -29 1415
rect -129 1365 -113 1399
rect -45 1365 -29 1399
rect -129 1318 -29 1365
rect 29 1399 129 1415
rect 29 1365 45 1399
rect 113 1365 129 1399
rect 29 1318 129 1365
rect 187 1399 287 1415
rect 187 1365 203 1399
rect 271 1365 287 1399
rect 187 1318 287 1365
rect 345 1399 445 1415
rect 345 1365 361 1399
rect 429 1365 445 1399
rect 345 1318 445 1365
rect 503 1399 603 1415
rect 503 1365 519 1399
rect 587 1365 603 1399
rect 503 1318 603 1365
rect 661 1399 761 1415
rect 661 1365 677 1399
rect 745 1365 761 1399
rect 661 1318 761 1365
rect 819 1399 919 1415
rect 819 1365 835 1399
rect 903 1365 919 1399
rect 819 1318 919 1365
rect 977 1399 1077 1415
rect 977 1365 993 1399
rect 1061 1365 1077 1399
rect 977 1318 1077 1365
rect -1077 71 -977 118
rect -1077 37 -1061 71
rect -993 37 -977 71
rect -1077 21 -977 37
rect -919 71 -819 118
rect -919 37 -903 71
rect -835 37 -819 71
rect -919 21 -819 37
rect -761 71 -661 118
rect -761 37 -745 71
rect -677 37 -661 71
rect -761 21 -661 37
rect -603 71 -503 118
rect -603 37 -587 71
rect -519 37 -503 71
rect -603 21 -503 37
rect -445 71 -345 118
rect -445 37 -429 71
rect -361 37 -345 71
rect -445 21 -345 37
rect -287 71 -187 118
rect -287 37 -271 71
rect -203 37 -187 71
rect -287 21 -187 37
rect -129 71 -29 118
rect -129 37 -113 71
rect -45 37 -29 71
rect -129 21 -29 37
rect 29 71 129 118
rect 29 37 45 71
rect 113 37 129 71
rect 29 21 129 37
rect 187 71 287 118
rect 187 37 203 71
rect 271 37 287 71
rect 187 21 287 37
rect 345 71 445 118
rect 345 37 361 71
rect 429 37 445 71
rect 345 21 445 37
rect 503 71 603 118
rect 503 37 519 71
rect 587 37 603 71
rect 503 21 603 37
rect 661 71 761 118
rect 661 37 677 71
rect 745 37 761 71
rect 661 21 761 37
rect 819 71 919 118
rect 819 37 835 71
rect 903 37 919 71
rect 819 21 919 37
rect 977 71 1077 118
rect 977 37 993 71
rect 1061 37 1077 71
rect 977 21 1077 37
rect -1077 -37 -977 -21
rect -1077 -71 -1061 -37
rect -993 -71 -977 -37
rect -1077 -118 -977 -71
rect -919 -37 -819 -21
rect -919 -71 -903 -37
rect -835 -71 -819 -37
rect -919 -118 -819 -71
rect -761 -37 -661 -21
rect -761 -71 -745 -37
rect -677 -71 -661 -37
rect -761 -118 -661 -71
rect -603 -37 -503 -21
rect -603 -71 -587 -37
rect -519 -71 -503 -37
rect -603 -118 -503 -71
rect -445 -37 -345 -21
rect -445 -71 -429 -37
rect -361 -71 -345 -37
rect -445 -118 -345 -71
rect -287 -37 -187 -21
rect -287 -71 -271 -37
rect -203 -71 -187 -37
rect -287 -118 -187 -71
rect -129 -37 -29 -21
rect -129 -71 -113 -37
rect -45 -71 -29 -37
rect -129 -118 -29 -71
rect 29 -37 129 -21
rect 29 -71 45 -37
rect 113 -71 129 -37
rect 29 -118 129 -71
rect 187 -37 287 -21
rect 187 -71 203 -37
rect 271 -71 287 -37
rect 187 -118 287 -71
rect 345 -37 445 -21
rect 345 -71 361 -37
rect 429 -71 445 -37
rect 345 -118 445 -71
rect 503 -37 603 -21
rect 503 -71 519 -37
rect 587 -71 603 -37
rect 503 -118 603 -71
rect 661 -37 761 -21
rect 661 -71 677 -37
rect 745 -71 761 -37
rect 661 -118 761 -71
rect 819 -37 919 -21
rect 819 -71 835 -37
rect 903 -71 919 -37
rect 819 -118 919 -71
rect 977 -37 1077 -21
rect 977 -71 993 -37
rect 1061 -71 1077 -37
rect 977 -118 1077 -71
rect -1077 -1365 -977 -1318
rect -1077 -1399 -1061 -1365
rect -993 -1399 -977 -1365
rect -1077 -1415 -977 -1399
rect -919 -1365 -819 -1318
rect -919 -1399 -903 -1365
rect -835 -1399 -819 -1365
rect -919 -1415 -819 -1399
rect -761 -1365 -661 -1318
rect -761 -1399 -745 -1365
rect -677 -1399 -661 -1365
rect -761 -1415 -661 -1399
rect -603 -1365 -503 -1318
rect -603 -1399 -587 -1365
rect -519 -1399 -503 -1365
rect -603 -1415 -503 -1399
rect -445 -1365 -345 -1318
rect -445 -1399 -429 -1365
rect -361 -1399 -345 -1365
rect -445 -1415 -345 -1399
rect -287 -1365 -187 -1318
rect -287 -1399 -271 -1365
rect -203 -1399 -187 -1365
rect -287 -1415 -187 -1399
rect -129 -1365 -29 -1318
rect -129 -1399 -113 -1365
rect -45 -1399 -29 -1365
rect -129 -1415 -29 -1399
rect 29 -1365 129 -1318
rect 29 -1399 45 -1365
rect 113 -1399 129 -1365
rect 29 -1415 129 -1399
rect 187 -1365 287 -1318
rect 187 -1399 203 -1365
rect 271 -1399 287 -1365
rect 187 -1415 287 -1399
rect 345 -1365 445 -1318
rect 345 -1399 361 -1365
rect 429 -1399 445 -1365
rect 345 -1415 445 -1399
rect 503 -1365 603 -1318
rect 503 -1399 519 -1365
rect 587 -1399 603 -1365
rect 503 -1415 603 -1399
rect 661 -1365 761 -1318
rect 661 -1399 677 -1365
rect 745 -1399 761 -1365
rect 661 -1415 761 -1399
rect 819 -1365 919 -1318
rect 819 -1399 835 -1365
rect 903 -1399 919 -1365
rect 819 -1415 919 -1399
rect 977 -1365 1077 -1318
rect 977 -1399 993 -1365
rect 1061 -1399 1077 -1365
rect 977 -1415 1077 -1399
rect -1077 -1473 -977 -1457
rect -1077 -1507 -1061 -1473
rect -993 -1507 -977 -1473
rect -1077 -1554 -977 -1507
rect -919 -1473 -819 -1457
rect -919 -1507 -903 -1473
rect -835 -1507 -819 -1473
rect -919 -1554 -819 -1507
rect -761 -1473 -661 -1457
rect -761 -1507 -745 -1473
rect -677 -1507 -661 -1473
rect -761 -1554 -661 -1507
rect -603 -1473 -503 -1457
rect -603 -1507 -587 -1473
rect -519 -1507 -503 -1473
rect -603 -1554 -503 -1507
rect -445 -1473 -345 -1457
rect -445 -1507 -429 -1473
rect -361 -1507 -345 -1473
rect -445 -1554 -345 -1507
rect -287 -1473 -187 -1457
rect -287 -1507 -271 -1473
rect -203 -1507 -187 -1473
rect -287 -1554 -187 -1507
rect -129 -1473 -29 -1457
rect -129 -1507 -113 -1473
rect -45 -1507 -29 -1473
rect -129 -1554 -29 -1507
rect 29 -1473 129 -1457
rect 29 -1507 45 -1473
rect 113 -1507 129 -1473
rect 29 -1554 129 -1507
rect 187 -1473 287 -1457
rect 187 -1507 203 -1473
rect 271 -1507 287 -1473
rect 187 -1554 287 -1507
rect 345 -1473 445 -1457
rect 345 -1507 361 -1473
rect 429 -1507 445 -1473
rect 345 -1554 445 -1507
rect 503 -1473 603 -1457
rect 503 -1507 519 -1473
rect 587 -1507 603 -1473
rect 503 -1554 603 -1507
rect 661 -1473 761 -1457
rect 661 -1507 677 -1473
rect 745 -1507 761 -1473
rect 661 -1554 761 -1507
rect 819 -1473 919 -1457
rect 819 -1507 835 -1473
rect 903 -1507 919 -1473
rect 819 -1554 919 -1507
rect 977 -1473 1077 -1457
rect 977 -1507 993 -1473
rect 1061 -1507 1077 -1473
rect 977 -1554 1077 -1507
rect -1077 -2801 -977 -2754
rect -1077 -2835 -1061 -2801
rect -993 -2835 -977 -2801
rect -1077 -2851 -977 -2835
rect -919 -2801 -819 -2754
rect -919 -2835 -903 -2801
rect -835 -2835 -819 -2801
rect -919 -2851 -819 -2835
rect -761 -2801 -661 -2754
rect -761 -2835 -745 -2801
rect -677 -2835 -661 -2801
rect -761 -2851 -661 -2835
rect -603 -2801 -503 -2754
rect -603 -2835 -587 -2801
rect -519 -2835 -503 -2801
rect -603 -2851 -503 -2835
rect -445 -2801 -345 -2754
rect -445 -2835 -429 -2801
rect -361 -2835 -345 -2801
rect -445 -2851 -345 -2835
rect -287 -2801 -187 -2754
rect -287 -2835 -271 -2801
rect -203 -2835 -187 -2801
rect -287 -2851 -187 -2835
rect -129 -2801 -29 -2754
rect -129 -2835 -113 -2801
rect -45 -2835 -29 -2801
rect -129 -2851 -29 -2835
rect 29 -2801 129 -2754
rect 29 -2835 45 -2801
rect 113 -2835 129 -2801
rect 29 -2851 129 -2835
rect 187 -2801 287 -2754
rect 187 -2835 203 -2801
rect 271 -2835 287 -2801
rect 187 -2851 287 -2835
rect 345 -2801 445 -2754
rect 345 -2835 361 -2801
rect 429 -2835 445 -2801
rect 345 -2851 445 -2835
rect 503 -2801 603 -2754
rect 503 -2835 519 -2801
rect 587 -2835 603 -2801
rect 503 -2851 603 -2835
rect 661 -2801 761 -2754
rect 661 -2835 677 -2801
rect 745 -2835 761 -2801
rect 661 -2851 761 -2835
rect 819 -2801 919 -2754
rect 819 -2835 835 -2801
rect 903 -2835 919 -2801
rect 819 -2851 919 -2835
rect 977 -2801 1077 -2754
rect 977 -2835 993 -2801
rect 1061 -2835 1077 -2801
rect 977 -2851 1077 -2835
<< polycont >>
rect -1061 2801 -993 2835
rect -903 2801 -835 2835
rect -745 2801 -677 2835
rect -587 2801 -519 2835
rect -429 2801 -361 2835
rect -271 2801 -203 2835
rect -113 2801 -45 2835
rect 45 2801 113 2835
rect 203 2801 271 2835
rect 361 2801 429 2835
rect 519 2801 587 2835
rect 677 2801 745 2835
rect 835 2801 903 2835
rect 993 2801 1061 2835
rect -1061 1473 -993 1507
rect -903 1473 -835 1507
rect -745 1473 -677 1507
rect -587 1473 -519 1507
rect -429 1473 -361 1507
rect -271 1473 -203 1507
rect -113 1473 -45 1507
rect 45 1473 113 1507
rect 203 1473 271 1507
rect 361 1473 429 1507
rect 519 1473 587 1507
rect 677 1473 745 1507
rect 835 1473 903 1507
rect 993 1473 1061 1507
rect -1061 1365 -993 1399
rect -903 1365 -835 1399
rect -745 1365 -677 1399
rect -587 1365 -519 1399
rect -429 1365 -361 1399
rect -271 1365 -203 1399
rect -113 1365 -45 1399
rect 45 1365 113 1399
rect 203 1365 271 1399
rect 361 1365 429 1399
rect 519 1365 587 1399
rect 677 1365 745 1399
rect 835 1365 903 1399
rect 993 1365 1061 1399
rect -1061 37 -993 71
rect -903 37 -835 71
rect -745 37 -677 71
rect -587 37 -519 71
rect -429 37 -361 71
rect -271 37 -203 71
rect -113 37 -45 71
rect 45 37 113 71
rect 203 37 271 71
rect 361 37 429 71
rect 519 37 587 71
rect 677 37 745 71
rect 835 37 903 71
rect 993 37 1061 71
rect -1061 -71 -993 -37
rect -903 -71 -835 -37
rect -745 -71 -677 -37
rect -587 -71 -519 -37
rect -429 -71 -361 -37
rect -271 -71 -203 -37
rect -113 -71 -45 -37
rect 45 -71 113 -37
rect 203 -71 271 -37
rect 361 -71 429 -37
rect 519 -71 587 -37
rect 677 -71 745 -37
rect 835 -71 903 -37
rect 993 -71 1061 -37
rect -1061 -1399 -993 -1365
rect -903 -1399 -835 -1365
rect -745 -1399 -677 -1365
rect -587 -1399 -519 -1365
rect -429 -1399 -361 -1365
rect -271 -1399 -203 -1365
rect -113 -1399 -45 -1365
rect 45 -1399 113 -1365
rect 203 -1399 271 -1365
rect 361 -1399 429 -1365
rect 519 -1399 587 -1365
rect 677 -1399 745 -1365
rect 835 -1399 903 -1365
rect 993 -1399 1061 -1365
rect -1061 -1507 -993 -1473
rect -903 -1507 -835 -1473
rect -745 -1507 -677 -1473
rect -587 -1507 -519 -1473
rect -429 -1507 -361 -1473
rect -271 -1507 -203 -1473
rect -113 -1507 -45 -1473
rect 45 -1507 113 -1473
rect 203 -1507 271 -1473
rect 361 -1507 429 -1473
rect 519 -1507 587 -1473
rect 677 -1507 745 -1473
rect 835 -1507 903 -1473
rect 993 -1507 1061 -1473
rect -1061 -2835 -993 -2801
rect -903 -2835 -835 -2801
rect -745 -2835 -677 -2801
rect -587 -2835 -519 -2801
rect -429 -2835 -361 -2801
rect -271 -2835 -203 -2801
rect -113 -2835 -45 -2801
rect 45 -2835 113 -2801
rect 203 -2835 271 -2801
rect 361 -2835 429 -2801
rect 519 -2835 587 -2801
rect 677 -2835 745 -2801
rect 835 -2835 903 -2801
rect 993 -2835 1061 -2801
<< locali >>
rect -1237 2903 -1141 2937
rect 1141 2903 1237 2937
rect -1237 2841 -1203 2903
rect 1203 2841 1237 2903
rect -1077 2801 -1061 2835
rect -993 2801 -977 2835
rect -919 2801 -903 2835
rect -835 2801 -819 2835
rect -761 2801 -745 2835
rect -677 2801 -661 2835
rect -603 2801 -587 2835
rect -519 2801 -503 2835
rect -445 2801 -429 2835
rect -361 2801 -345 2835
rect -287 2801 -271 2835
rect -203 2801 -187 2835
rect -129 2801 -113 2835
rect -45 2801 -29 2835
rect 29 2801 45 2835
rect 113 2801 129 2835
rect 187 2801 203 2835
rect 271 2801 287 2835
rect 345 2801 361 2835
rect 429 2801 445 2835
rect 503 2801 519 2835
rect 587 2801 603 2835
rect 661 2801 677 2835
rect 745 2801 761 2835
rect 819 2801 835 2835
rect 903 2801 919 2835
rect 977 2801 993 2835
rect 1061 2801 1077 2835
rect -1123 2742 -1089 2758
rect -1123 1550 -1089 1566
rect -965 2742 -931 2758
rect -965 1550 -931 1566
rect -807 2742 -773 2758
rect -807 1550 -773 1566
rect -649 2742 -615 2758
rect -649 1550 -615 1566
rect -491 2742 -457 2758
rect -491 1550 -457 1566
rect -333 2742 -299 2758
rect -333 1550 -299 1566
rect -175 2742 -141 2758
rect -175 1550 -141 1566
rect -17 2742 17 2758
rect -17 1550 17 1566
rect 141 2742 175 2758
rect 141 1550 175 1566
rect 299 2742 333 2758
rect 299 1550 333 1566
rect 457 2742 491 2758
rect 457 1550 491 1566
rect 615 2742 649 2758
rect 615 1550 649 1566
rect 773 2742 807 2758
rect 773 1550 807 1566
rect 931 2742 965 2758
rect 931 1550 965 1566
rect 1089 2742 1123 2758
rect 1089 1550 1123 1566
rect -1077 1473 -1061 1507
rect -993 1473 -977 1507
rect -919 1473 -903 1507
rect -835 1473 -819 1507
rect -761 1473 -745 1507
rect -677 1473 -661 1507
rect -603 1473 -587 1507
rect -519 1473 -503 1507
rect -445 1473 -429 1507
rect -361 1473 -345 1507
rect -287 1473 -271 1507
rect -203 1473 -187 1507
rect -129 1473 -113 1507
rect -45 1473 -29 1507
rect 29 1473 45 1507
rect 113 1473 129 1507
rect 187 1473 203 1507
rect 271 1473 287 1507
rect 345 1473 361 1507
rect 429 1473 445 1507
rect 503 1473 519 1507
rect 587 1473 603 1507
rect 661 1473 677 1507
rect 745 1473 761 1507
rect 819 1473 835 1507
rect 903 1473 919 1507
rect 977 1473 993 1507
rect 1061 1473 1077 1507
rect -1077 1365 -1061 1399
rect -993 1365 -977 1399
rect -919 1365 -903 1399
rect -835 1365 -819 1399
rect -761 1365 -745 1399
rect -677 1365 -661 1399
rect -603 1365 -587 1399
rect -519 1365 -503 1399
rect -445 1365 -429 1399
rect -361 1365 -345 1399
rect -287 1365 -271 1399
rect -203 1365 -187 1399
rect -129 1365 -113 1399
rect -45 1365 -29 1399
rect 29 1365 45 1399
rect 113 1365 129 1399
rect 187 1365 203 1399
rect 271 1365 287 1399
rect 345 1365 361 1399
rect 429 1365 445 1399
rect 503 1365 519 1399
rect 587 1365 603 1399
rect 661 1365 677 1399
rect 745 1365 761 1399
rect 819 1365 835 1399
rect 903 1365 919 1399
rect 977 1365 993 1399
rect 1061 1365 1077 1399
rect -1123 1306 -1089 1322
rect -1123 114 -1089 130
rect -965 1306 -931 1322
rect -965 114 -931 130
rect -807 1306 -773 1322
rect -807 114 -773 130
rect -649 1306 -615 1322
rect -649 114 -615 130
rect -491 1306 -457 1322
rect -491 114 -457 130
rect -333 1306 -299 1322
rect -333 114 -299 130
rect -175 1306 -141 1322
rect -175 114 -141 130
rect -17 1306 17 1322
rect -17 114 17 130
rect 141 1306 175 1322
rect 141 114 175 130
rect 299 1306 333 1322
rect 299 114 333 130
rect 457 1306 491 1322
rect 457 114 491 130
rect 615 1306 649 1322
rect 615 114 649 130
rect 773 1306 807 1322
rect 773 114 807 130
rect 931 1306 965 1322
rect 931 114 965 130
rect 1089 1306 1123 1322
rect 1089 114 1123 130
rect -1077 37 -1061 71
rect -993 37 -977 71
rect -919 37 -903 71
rect -835 37 -819 71
rect -761 37 -745 71
rect -677 37 -661 71
rect -603 37 -587 71
rect -519 37 -503 71
rect -445 37 -429 71
rect -361 37 -345 71
rect -287 37 -271 71
rect -203 37 -187 71
rect -129 37 -113 71
rect -45 37 -29 71
rect 29 37 45 71
rect 113 37 129 71
rect 187 37 203 71
rect 271 37 287 71
rect 345 37 361 71
rect 429 37 445 71
rect 503 37 519 71
rect 587 37 603 71
rect 661 37 677 71
rect 745 37 761 71
rect 819 37 835 71
rect 903 37 919 71
rect 977 37 993 71
rect 1061 37 1077 71
rect -1077 -71 -1061 -37
rect -993 -71 -977 -37
rect -919 -71 -903 -37
rect -835 -71 -819 -37
rect -761 -71 -745 -37
rect -677 -71 -661 -37
rect -603 -71 -587 -37
rect -519 -71 -503 -37
rect -445 -71 -429 -37
rect -361 -71 -345 -37
rect -287 -71 -271 -37
rect -203 -71 -187 -37
rect -129 -71 -113 -37
rect -45 -71 -29 -37
rect 29 -71 45 -37
rect 113 -71 129 -37
rect 187 -71 203 -37
rect 271 -71 287 -37
rect 345 -71 361 -37
rect 429 -71 445 -37
rect 503 -71 519 -37
rect 587 -71 603 -37
rect 661 -71 677 -37
rect 745 -71 761 -37
rect 819 -71 835 -37
rect 903 -71 919 -37
rect 977 -71 993 -37
rect 1061 -71 1077 -37
rect -1123 -130 -1089 -114
rect -1123 -1322 -1089 -1306
rect -965 -130 -931 -114
rect -965 -1322 -931 -1306
rect -807 -130 -773 -114
rect -807 -1322 -773 -1306
rect -649 -130 -615 -114
rect -649 -1322 -615 -1306
rect -491 -130 -457 -114
rect -491 -1322 -457 -1306
rect -333 -130 -299 -114
rect -333 -1322 -299 -1306
rect -175 -130 -141 -114
rect -175 -1322 -141 -1306
rect -17 -130 17 -114
rect -17 -1322 17 -1306
rect 141 -130 175 -114
rect 141 -1322 175 -1306
rect 299 -130 333 -114
rect 299 -1322 333 -1306
rect 457 -130 491 -114
rect 457 -1322 491 -1306
rect 615 -130 649 -114
rect 615 -1322 649 -1306
rect 773 -130 807 -114
rect 773 -1322 807 -1306
rect 931 -130 965 -114
rect 931 -1322 965 -1306
rect 1089 -130 1123 -114
rect 1089 -1322 1123 -1306
rect -1077 -1399 -1061 -1365
rect -993 -1399 -977 -1365
rect -919 -1399 -903 -1365
rect -835 -1399 -819 -1365
rect -761 -1399 -745 -1365
rect -677 -1399 -661 -1365
rect -603 -1399 -587 -1365
rect -519 -1399 -503 -1365
rect -445 -1399 -429 -1365
rect -361 -1399 -345 -1365
rect -287 -1399 -271 -1365
rect -203 -1399 -187 -1365
rect -129 -1399 -113 -1365
rect -45 -1399 -29 -1365
rect 29 -1399 45 -1365
rect 113 -1399 129 -1365
rect 187 -1399 203 -1365
rect 271 -1399 287 -1365
rect 345 -1399 361 -1365
rect 429 -1399 445 -1365
rect 503 -1399 519 -1365
rect 587 -1399 603 -1365
rect 661 -1399 677 -1365
rect 745 -1399 761 -1365
rect 819 -1399 835 -1365
rect 903 -1399 919 -1365
rect 977 -1399 993 -1365
rect 1061 -1399 1077 -1365
rect -1077 -1507 -1061 -1473
rect -993 -1507 -977 -1473
rect -919 -1507 -903 -1473
rect -835 -1507 -819 -1473
rect -761 -1507 -745 -1473
rect -677 -1507 -661 -1473
rect -603 -1507 -587 -1473
rect -519 -1507 -503 -1473
rect -445 -1507 -429 -1473
rect -361 -1507 -345 -1473
rect -287 -1507 -271 -1473
rect -203 -1507 -187 -1473
rect -129 -1507 -113 -1473
rect -45 -1507 -29 -1473
rect 29 -1507 45 -1473
rect 113 -1507 129 -1473
rect 187 -1507 203 -1473
rect 271 -1507 287 -1473
rect 345 -1507 361 -1473
rect 429 -1507 445 -1473
rect 503 -1507 519 -1473
rect 587 -1507 603 -1473
rect 661 -1507 677 -1473
rect 745 -1507 761 -1473
rect 819 -1507 835 -1473
rect 903 -1507 919 -1473
rect 977 -1507 993 -1473
rect 1061 -1507 1077 -1473
rect -1123 -1566 -1089 -1550
rect -1123 -2758 -1089 -2742
rect -965 -1566 -931 -1550
rect -965 -2758 -931 -2742
rect -807 -1566 -773 -1550
rect -807 -2758 -773 -2742
rect -649 -1566 -615 -1550
rect -649 -2758 -615 -2742
rect -491 -1566 -457 -1550
rect -491 -2758 -457 -2742
rect -333 -1566 -299 -1550
rect -333 -2758 -299 -2742
rect -175 -1566 -141 -1550
rect -175 -2758 -141 -2742
rect -17 -1566 17 -1550
rect -17 -2758 17 -2742
rect 141 -1566 175 -1550
rect 141 -2758 175 -2742
rect 299 -1566 333 -1550
rect 299 -2758 333 -2742
rect 457 -1566 491 -1550
rect 457 -2758 491 -2742
rect 615 -1566 649 -1550
rect 615 -2758 649 -2742
rect 773 -1566 807 -1550
rect 773 -2758 807 -2742
rect 931 -1566 965 -1550
rect 931 -2758 965 -2742
rect 1089 -1566 1123 -1550
rect 1089 -2758 1123 -2742
rect -1077 -2835 -1061 -2801
rect -993 -2835 -977 -2801
rect -919 -2835 -903 -2801
rect -835 -2835 -819 -2801
rect -761 -2835 -745 -2801
rect -677 -2835 -661 -2801
rect -603 -2835 -587 -2801
rect -519 -2835 -503 -2801
rect -445 -2835 -429 -2801
rect -361 -2835 -345 -2801
rect -287 -2835 -271 -2801
rect -203 -2835 -187 -2801
rect -129 -2835 -113 -2801
rect -45 -2835 -29 -2801
rect 29 -2835 45 -2801
rect 113 -2835 129 -2801
rect 187 -2835 203 -2801
rect 271 -2835 287 -2801
rect 345 -2835 361 -2801
rect 429 -2835 445 -2801
rect 503 -2835 519 -2801
rect 587 -2835 603 -2801
rect 661 -2835 677 -2801
rect 745 -2835 761 -2801
rect 819 -2835 835 -2801
rect 903 -2835 919 -2801
rect 977 -2835 993 -2801
rect 1061 -2835 1077 -2801
rect -1237 -2903 -1203 -2841
rect 1203 -2903 1237 -2841
rect -1237 -2937 -1141 -2903
rect 1141 -2937 1237 -2903
<< viali >>
rect -1061 2801 -993 2835
rect -903 2801 -835 2835
rect -745 2801 -677 2835
rect -587 2801 -519 2835
rect -429 2801 -361 2835
rect -271 2801 -203 2835
rect -113 2801 -45 2835
rect 45 2801 113 2835
rect 203 2801 271 2835
rect 361 2801 429 2835
rect 519 2801 587 2835
rect 677 2801 745 2835
rect 835 2801 903 2835
rect 993 2801 1061 2835
rect -1123 1566 -1089 2742
rect -965 1566 -931 2742
rect -807 1566 -773 2742
rect -649 1566 -615 2742
rect -491 1566 -457 2742
rect -333 1566 -299 2742
rect -175 1566 -141 2742
rect -17 1566 17 2742
rect 141 1566 175 2742
rect 299 1566 333 2742
rect 457 1566 491 2742
rect 615 1566 649 2742
rect 773 1566 807 2742
rect 931 1566 965 2742
rect 1089 1566 1123 2742
rect -1061 1473 -993 1507
rect -903 1473 -835 1507
rect -745 1473 -677 1507
rect -587 1473 -519 1507
rect -429 1473 -361 1507
rect -271 1473 -203 1507
rect -113 1473 -45 1507
rect 45 1473 113 1507
rect 203 1473 271 1507
rect 361 1473 429 1507
rect 519 1473 587 1507
rect 677 1473 745 1507
rect 835 1473 903 1507
rect 993 1473 1061 1507
rect -1061 1365 -993 1399
rect -903 1365 -835 1399
rect -745 1365 -677 1399
rect -587 1365 -519 1399
rect -429 1365 -361 1399
rect -271 1365 -203 1399
rect -113 1365 -45 1399
rect 45 1365 113 1399
rect 203 1365 271 1399
rect 361 1365 429 1399
rect 519 1365 587 1399
rect 677 1365 745 1399
rect 835 1365 903 1399
rect 993 1365 1061 1399
rect -1123 130 -1089 1306
rect -965 130 -931 1306
rect -807 130 -773 1306
rect -649 130 -615 1306
rect -491 130 -457 1306
rect -333 130 -299 1306
rect -175 130 -141 1306
rect -17 130 17 1306
rect 141 130 175 1306
rect 299 130 333 1306
rect 457 130 491 1306
rect 615 130 649 1306
rect 773 130 807 1306
rect 931 130 965 1306
rect 1089 130 1123 1306
rect -1061 37 -993 71
rect -903 37 -835 71
rect -745 37 -677 71
rect -587 37 -519 71
rect -429 37 -361 71
rect -271 37 -203 71
rect -113 37 -45 71
rect 45 37 113 71
rect 203 37 271 71
rect 361 37 429 71
rect 519 37 587 71
rect 677 37 745 71
rect 835 37 903 71
rect 993 37 1061 71
rect -1061 -71 -993 -37
rect -903 -71 -835 -37
rect -745 -71 -677 -37
rect -587 -71 -519 -37
rect -429 -71 -361 -37
rect -271 -71 -203 -37
rect -113 -71 -45 -37
rect 45 -71 113 -37
rect 203 -71 271 -37
rect 361 -71 429 -37
rect 519 -71 587 -37
rect 677 -71 745 -37
rect 835 -71 903 -37
rect 993 -71 1061 -37
rect -1123 -1306 -1089 -130
rect -965 -1306 -931 -130
rect -807 -1306 -773 -130
rect -649 -1306 -615 -130
rect -491 -1306 -457 -130
rect -333 -1306 -299 -130
rect -175 -1306 -141 -130
rect -17 -1306 17 -130
rect 141 -1306 175 -130
rect 299 -1306 333 -130
rect 457 -1306 491 -130
rect 615 -1306 649 -130
rect 773 -1306 807 -130
rect 931 -1306 965 -130
rect 1089 -1306 1123 -130
rect -1061 -1399 -993 -1365
rect -903 -1399 -835 -1365
rect -745 -1399 -677 -1365
rect -587 -1399 -519 -1365
rect -429 -1399 -361 -1365
rect -271 -1399 -203 -1365
rect -113 -1399 -45 -1365
rect 45 -1399 113 -1365
rect 203 -1399 271 -1365
rect 361 -1399 429 -1365
rect 519 -1399 587 -1365
rect 677 -1399 745 -1365
rect 835 -1399 903 -1365
rect 993 -1399 1061 -1365
rect -1061 -1507 -993 -1473
rect -903 -1507 -835 -1473
rect -745 -1507 -677 -1473
rect -587 -1507 -519 -1473
rect -429 -1507 -361 -1473
rect -271 -1507 -203 -1473
rect -113 -1507 -45 -1473
rect 45 -1507 113 -1473
rect 203 -1507 271 -1473
rect 361 -1507 429 -1473
rect 519 -1507 587 -1473
rect 677 -1507 745 -1473
rect 835 -1507 903 -1473
rect 993 -1507 1061 -1473
rect -1123 -2742 -1089 -1566
rect -965 -2742 -931 -1566
rect -807 -2742 -773 -1566
rect -649 -2742 -615 -1566
rect -491 -2742 -457 -1566
rect -333 -2742 -299 -1566
rect -175 -2742 -141 -1566
rect -17 -2742 17 -1566
rect 141 -2742 175 -1566
rect 299 -2742 333 -1566
rect 457 -2742 491 -1566
rect 615 -2742 649 -1566
rect 773 -2742 807 -1566
rect 931 -2742 965 -1566
rect 1089 -2742 1123 -1566
rect -1061 -2835 -993 -2801
rect -903 -2835 -835 -2801
rect -745 -2835 -677 -2801
rect -587 -2835 -519 -2801
rect -429 -2835 -361 -2801
rect -271 -2835 -203 -2801
rect -113 -2835 -45 -2801
rect 45 -2835 113 -2801
rect 203 -2835 271 -2801
rect 361 -2835 429 -2801
rect 519 -2835 587 -2801
rect 677 -2835 745 -2801
rect 835 -2835 903 -2801
rect 993 -2835 1061 -2801
<< metal1 >>
rect -1073 2835 -981 2841
rect -1073 2801 -1061 2835
rect -993 2801 -981 2835
rect -1073 2795 -981 2801
rect -915 2835 -823 2841
rect -915 2801 -903 2835
rect -835 2801 -823 2835
rect -915 2795 -823 2801
rect -757 2835 -665 2841
rect -757 2801 -745 2835
rect -677 2801 -665 2835
rect -757 2795 -665 2801
rect -599 2835 -507 2841
rect -599 2801 -587 2835
rect -519 2801 -507 2835
rect -599 2795 -507 2801
rect -441 2835 -349 2841
rect -441 2801 -429 2835
rect -361 2801 -349 2835
rect -441 2795 -349 2801
rect -283 2835 -191 2841
rect -283 2801 -271 2835
rect -203 2801 -191 2835
rect -283 2795 -191 2801
rect -125 2835 -33 2841
rect -125 2801 -113 2835
rect -45 2801 -33 2835
rect -125 2795 -33 2801
rect 33 2835 125 2841
rect 33 2801 45 2835
rect 113 2801 125 2835
rect 33 2795 125 2801
rect 191 2835 283 2841
rect 191 2801 203 2835
rect 271 2801 283 2835
rect 191 2795 283 2801
rect 349 2835 441 2841
rect 349 2801 361 2835
rect 429 2801 441 2835
rect 349 2795 441 2801
rect 507 2835 599 2841
rect 507 2801 519 2835
rect 587 2801 599 2835
rect 507 2795 599 2801
rect 665 2835 757 2841
rect 665 2801 677 2835
rect 745 2801 757 2835
rect 665 2795 757 2801
rect 823 2835 915 2841
rect 823 2801 835 2835
rect 903 2801 915 2835
rect 823 2795 915 2801
rect 981 2835 1073 2841
rect 981 2801 993 2835
rect 1061 2801 1073 2835
rect 981 2795 1073 2801
rect -1129 2742 -1083 2754
rect -1129 1566 -1123 2742
rect -1089 1566 -1083 2742
rect -1129 1554 -1083 1566
rect -971 2742 -925 2754
rect -971 1566 -965 2742
rect -931 1566 -925 2742
rect -971 1554 -925 1566
rect -813 2742 -767 2754
rect -813 1566 -807 2742
rect -773 1566 -767 2742
rect -813 1554 -767 1566
rect -655 2742 -609 2754
rect -655 1566 -649 2742
rect -615 1566 -609 2742
rect -655 1554 -609 1566
rect -497 2742 -451 2754
rect -497 1566 -491 2742
rect -457 1566 -451 2742
rect -497 1554 -451 1566
rect -339 2742 -293 2754
rect -339 1566 -333 2742
rect -299 1566 -293 2742
rect -339 1554 -293 1566
rect -181 2742 -135 2754
rect -181 1566 -175 2742
rect -141 1566 -135 2742
rect -181 1554 -135 1566
rect -23 2742 23 2754
rect -23 1566 -17 2742
rect 17 1566 23 2742
rect -23 1554 23 1566
rect 135 2742 181 2754
rect 135 1566 141 2742
rect 175 1566 181 2742
rect 135 1554 181 1566
rect 293 2742 339 2754
rect 293 1566 299 2742
rect 333 1566 339 2742
rect 293 1554 339 1566
rect 451 2742 497 2754
rect 451 1566 457 2742
rect 491 1566 497 2742
rect 451 1554 497 1566
rect 609 2742 655 2754
rect 609 1566 615 2742
rect 649 1566 655 2742
rect 609 1554 655 1566
rect 767 2742 813 2754
rect 767 1566 773 2742
rect 807 1566 813 2742
rect 767 1554 813 1566
rect 925 2742 971 2754
rect 925 1566 931 2742
rect 965 1566 971 2742
rect 925 1554 971 1566
rect 1083 2742 1129 2754
rect 1083 1566 1089 2742
rect 1123 1566 1129 2742
rect 1083 1554 1129 1566
rect -1073 1507 -981 1513
rect -1073 1473 -1061 1507
rect -993 1473 -981 1507
rect -1073 1467 -981 1473
rect -915 1507 -823 1513
rect -915 1473 -903 1507
rect -835 1473 -823 1507
rect -915 1467 -823 1473
rect -757 1507 -665 1513
rect -757 1473 -745 1507
rect -677 1473 -665 1507
rect -757 1467 -665 1473
rect -599 1507 -507 1513
rect -599 1473 -587 1507
rect -519 1473 -507 1507
rect -599 1467 -507 1473
rect -441 1507 -349 1513
rect -441 1473 -429 1507
rect -361 1473 -349 1507
rect -441 1467 -349 1473
rect -283 1507 -191 1513
rect -283 1473 -271 1507
rect -203 1473 -191 1507
rect -283 1467 -191 1473
rect -125 1507 -33 1513
rect -125 1473 -113 1507
rect -45 1473 -33 1507
rect -125 1467 -33 1473
rect 33 1507 125 1513
rect 33 1473 45 1507
rect 113 1473 125 1507
rect 33 1467 125 1473
rect 191 1507 283 1513
rect 191 1473 203 1507
rect 271 1473 283 1507
rect 191 1467 283 1473
rect 349 1507 441 1513
rect 349 1473 361 1507
rect 429 1473 441 1507
rect 349 1467 441 1473
rect 507 1507 599 1513
rect 507 1473 519 1507
rect 587 1473 599 1507
rect 507 1467 599 1473
rect 665 1507 757 1513
rect 665 1473 677 1507
rect 745 1473 757 1507
rect 665 1467 757 1473
rect 823 1507 915 1513
rect 823 1473 835 1507
rect 903 1473 915 1507
rect 823 1467 915 1473
rect 981 1507 1073 1513
rect 981 1473 993 1507
rect 1061 1473 1073 1507
rect 981 1467 1073 1473
rect -1073 1399 -981 1405
rect -1073 1365 -1061 1399
rect -993 1365 -981 1399
rect -1073 1359 -981 1365
rect -915 1399 -823 1405
rect -915 1365 -903 1399
rect -835 1365 -823 1399
rect -915 1359 -823 1365
rect -757 1399 -665 1405
rect -757 1365 -745 1399
rect -677 1365 -665 1399
rect -757 1359 -665 1365
rect -599 1399 -507 1405
rect -599 1365 -587 1399
rect -519 1365 -507 1399
rect -599 1359 -507 1365
rect -441 1399 -349 1405
rect -441 1365 -429 1399
rect -361 1365 -349 1399
rect -441 1359 -349 1365
rect -283 1399 -191 1405
rect -283 1365 -271 1399
rect -203 1365 -191 1399
rect -283 1359 -191 1365
rect -125 1399 -33 1405
rect -125 1365 -113 1399
rect -45 1365 -33 1399
rect -125 1359 -33 1365
rect 33 1399 125 1405
rect 33 1365 45 1399
rect 113 1365 125 1399
rect 33 1359 125 1365
rect 191 1399 283 1405
rect 191 1365 203 1399
rect 271 1365 283 1399
rect 191 1359 283 1365
rect 349 1399 441 1405
rect 349 1365 361 1399
rect 429 1365 441 1399
rect 349 1359 441 1365
rect 507 1399 599 1405
rect 507 1365 519 1399
rect 587 1365 599 1399
rect 507 1359 599 1365
rect 665 1399 757 1405
rect 665 1365 677 1399
rect 745 1365 757 1399
rect 665 1359 757 1365
rect 823 1399 915 1405
rect 823 1365 835 1399
rect 903 1365 915 1399
rect 823 1359 915 1365
rect 981 1399 1073 1405
rect 981 1365 993 1399
rect 1061 1365 1073 1399
rect 981 1359 1073 1365
rect -1129 1306 -1083 1318
rect -1129 130 -1123 1306
rect -1089 130 -1083 1306
rect -1129 118 -1083 130
rect -971 1306 -925 1318
rect -971 130 -965 1306
rect -931 130 -925 1306
rect -971 118 -925 130
rect -813 1306 -767 1318
rect -813 130 -807 1306
rect -773 130 -767 1306
rect -813 118 -767 130
rect -655 1306 -609 1318
rect -655 130 -649 1306
rect -615 130 -609 1306
rect -655 118 -609 130
rect -497 1306 -451 1318
rect -497 130 -491 1306
rect -457 130 -451 1306
rect -497 118 -451 130
rect -339 1306 -293 1318
rect -339 130 -333 1306
rect -299 130 -293 1306
rect -339 118 -293 130
rect -181 1306 -135 1318
rect -181 130 -175 1306
rect -141 130 -135 1306
rect -181 118 -135 130
rect -23 1306 23 1318
rect -23 130 -17 1306
rect 17 130 23 1306
rect -23 118 23 130
rect 135 1306 181 1318
rect 135 130 141 1306
rect 175 130 181 1306
rect 135 118 181 130
rect 293 1306 339 1318
rect 293 130 299 1306
rect 333 130 339 1306
rect 293 118 339 130
rect 451 1306 497 1318
rect 451 130 457 1306
rect 491 130 497 1306
rect 451 118 497 130
rect 609 1306 655 1318
rect 609 130 615 1306
rect 649 130 655 1306
rect 609 118 655 130
rect 767 1306 813 1318
rect 767 130 773 1306
rect 807 130 813 1306
rect 767 118 813 130
rect 925 1306 971 1318
rect 925 130 931 1306
rect 965 130 971 1306
rect 925 118 971 130
rect 1083 1306 1129 1318
rect 1083 130 1089 1306
rect 1123 130 1129 1306
rect 1083 118 1129 130
rect -1073 71 -981 77
rect -1073 37 -1061 71
rect -993 37 -981 71
rect -1073 31 -981 37
rect -915 71 -823 77
rect -915 37 -903 71
rect -835 37 -823 71
rect -915 31 -823 37
rect -757 71 -665 77
rect -757 37 -745 71
rect -677 37 -665 71
rect -757 31 -665 37
rect -599 71 -507 77
rect -599 37 -587 71
rect -519 37 -507 71
rect -599 31 -507 37
rect -441 71 -349 77
rect -441 37 -429 71
rect -361 37 -349 71
rect -441 31 -349 37
rect -283 71 -191 77
rect -283 37 -271 71
rect -203 37 -191 71
rect -283 31 -191 37
rect -125 71 -33 77
rect -125 37 -113 71
rect -45 37 -33 71
rect -125 31 -33 37
rect 33 71 125 77
rect 33 37 45 71
rect 113 37 125 71
rect 33 31 125 37
rect 191 71 283 77
rect 191 37 203 71
rect 271 37 283 71
rect 191 31 283 37
rect 349 71 441 77
rect 349 37 361 71
rect 429 37 441 71
rect 349 31 441 37
rect 507 71 599 77
rect 507 37 519 71
rect 587 37 599 71
rect 507 31 599 37
rect 665 71 757 77
rect 665 37 677 71
rect 745 37 757 71
rect 665 31 757 37
rect 823 71 915 77
rect 823 37 835 71
rect 903 37 915 71
rect 823 31 915 37
rect 981 71 1073 77
rect 981 37 993 71
rect 1061 37 1073 71
rect 981 31 1073 37
rect -1073 -37 -981 -31
rect -1073 -71 -1061 -37
rect -993 -71 -981 -37
rect -1073 -77 -981 -71
rect -915 -37 -823 -31
rect -915 -71 -903 -37
rect -835 -71 -823 -37
rect -915 -77 -823 -71
rect -757 -37 -665 -31
rect -757 -71 -745 -37
rect -677 -71 -665 -37
rect -757 -77 -665 -71
rect -599 -37 -507 -31
rect -599 -71 -587 -37
rect -519 -71 -507 -37
rect -599 -77 -507 -71
rect -441 -37 -349 -31
rect -441 -71 -429 -37
rect -361 -71 -349 -37
rect -441 -77 -349 -71
rect -283 -37 -191 -31
rect -283 -71 -271 -37
rect -203 -71 -191 -37
rect -283 -77 -191 -71
rect -125 -37 -33 -31
rect -125 -71 -113 -37
rect -45 -71 -33 -37
rect -125 -77 -33 -71
rect 33 -37 125 -31
rect 33 -71 45 -37
rect 113 -71 125 -37
rect 33 -77 125 -71
rect 191 -37 283 -31
rect 191 -71 203 -37
rect 271 -71 283 -37
rect 191 -77 283 -71
rect 349 -37 441 -31
rect 349 -71 361 -37
rect 429 -71 441 -37
rect 349 -77 441 -71
rect 507 -37 599 -31
rect 507 -71 519 -37
rect 587 -71 599 -37
rect 507 -77 599 -71
rect 665 -37 757 -31
rect 665 -71 677 -37
rect 745 -71 757 -37
rect 665 -77 757 -71
rect 823 -37 915 -31
rect 823 -71 835 -37
rect 903 -71 915 -37
rect 823 -77 915 -71
rect 981 -37 1073 -31
rect 981 -71 993 -37
rect 1061 -71 1073 -37
rect 981 -77 1073 -71
rect -1129 -130 -1083 -118
rect -1129 -1306 -1123 -130
rect -1089 -1306 -1083 -130
rect -1129 -1318 -1083 -1306
rect -971 -130 -925 -118
rect -971 -1306 -965 -130
rect -931 -1306 -925 -130
rect -971 -1318 -925 -1306
rect -813 -130 -767 -118
rect -813 -1306 -807 -130
rect -773 -1306 -767 -130
rect -813 -1318 -767 -1306
rect -655 -130 -609 -118
rect -655 -1306 -649 -130
rect -615 -1306 -609 -130
rect -655 -1318 -609 -1306
rect -497 -130 -451 -118
rect -497 -1306 -491 -130
rect -457 -1306 -451 -130
rect -497 -1318 -451 -1306
rect -339 -130 -293 -118
rect -339 -1306 -333 -130
rect -299 -1306 -293 -130
rect -339 -1318 -293 -1306
rect -181 -130 -135 -118
rect -181 -1306 -175 -130
rect -141 -1306 -135 -130
rect -181 -1318 -135 -1306
rect -23 -130 23 -118
rect -23 -1306 -17 -130
rect 17 -1306 23 -130
rect -23 -1318 23 -1306
rect 135 -130 181 -118
rect 135 -1306 141 -130
rect 175 -1306 181 -130
rect 135 -1318 181 -1306
rect 293 -130 339 -118
rect 293 -1306 299 -130
rect 333 -1306 339 -130
rect 293 -1318 339 -1306
rect 451 -130 497 -118
rect 451 -1306 457 -130
rect 491 -1306 497 -130
rect 451 -1318 497 -1306
rect 609 -130 655 -118
rect 609 -1306 615 -130
rect 649 -1306 655 -130
rect 609 -1318 655 -1306
rect 767 -130 813 -118
rect 767 -1306 773 -130
rect 807 -1306 813 -130
rect 767 -1318 813 -1306
rect 925 -130 971 -118
rect 925 -1306 931 -130
rect 965 -1306 971 -130
rect 925 -1318 971 -1306
rect 1083 -130 1129 -118
rect 1083 -1306 1089 -130
rect 1123 -1306 1129 -130
rect 1083 -1318 1129 -1306
rect -1073 -1365 -981 -1359
rect -1073 -1399 -1061 -1365
rect -993 -1399 -981 -1365
rect -1073 -1405 -981 -1399
rect -915 -1365 -823 -1359
rect -915 -1399 -903 -1365
rect -835 -1399 -823 -1365
rect -915 -1405 -823 -1399
rect -757 -1365 -665 -1359
rect -757 -1399 -745 -1365
rect -677 -1399 -665 -1365
rect -757 -1405 -665 -1399
rect -599 -1365 -507 -1359
rect -599 -1399 -587 -1365
rect -519 -1399 -507 -1365
rect -599 -1405 -507 -1399
rect -441 -1365 -349 -1359
rect -441 -1399 -429 -1365
rect -361 -1399 -349 -1365
rect -441 -1405 -349 -1399
rect -283 -1365 -191 -1359
rect -283 -1399 -271 -1365
rect -203 -1399 -191 -1365
rect -283 -1405 -191 -1399
rect -125 -1365 -33 -1359
rect -125 -1399 -113 -1365
rect -45 -1399 -33 -1365
rect -125 -1405 -33 -1399
rect 33 -1365 125 -1359
rect 33 -1399 45 -1365
rect 113 -1399 125 -1365
rect 33 -1405 125 -1399
rect 191 -1365 283 -1359
rect 191 -1399 203 -1365
rect 271 -1399 283 -1365
rect 191 -1405 283 -1399
rect 349 -1365 441 -1359
rect 349 -1399 361 -1365
rect 429 -1399 441 -1365
rect 349 -1405 441 -1399
rect 507 -1365 599 -1359
rect 507 -1399 519 -1365
rect 587 -1399 599 -1365
rect 507 -1405 599 -1399
rect 665 -1365 757 -1359
rect 665 -1399 677 -1365
rect 745 -1399 757 -1365
rect 665 -1405 757 -1399
rect 823 -1365 915 -1359
rect 823 -1399 835 -1365
rect 903 -1399 915 -1365
rect 823 -1405 915 -1399
rect 981 -1365 1073 -1359
rect 981 -1399 993 -1365
rect 1061 -1399 1073 -1365
rect 981 -1405 1073 -1399
rect -1073 -1473 -981 -1467
rect -1073 -1507 -1061 -1473
rect -993 -1507 -981 -1473
rect -1073 -1513 -981 -1507
rect -915 -1473 -823 -1467
rect -915 -1507 -903 -1473
rect -835 -1507 -823 -1473
rect -915 -1513 -823 -1507
rect -757 -1473 -665 -1467
rect -757 -1507 -745 -1473
rect -677 -1507 -665 -1473
rect -757 -1513 -665 -1507
rect -599 -1473 -507 -1467
rect -599 -1507 -587 -1473
rect -519 -1507 -507 -1473
rect -599 -1513 -507 -1507
rect -441 -1473 -349 -1467
rect -441 -1507 -429 -1473
rect -361 -1507 -349 -1473
rect -441 -1513 -349 -1507
rect -283 -1473 -191 -1467
rect -283 -1507 -271 -1473
rect -203 -1507 -191 -1473
rect -283 -1513 -191 -1507
rect -125 -1473 -33 -1467
rect -125 -1507 -113 -1473
rect -45 -1507 -33 -1473
rect -125 -1513 -33 -1507
rect 33 -1473 125 -1467
rect 33 -1507 45 -1473
rect 113 -1507 125 -1473
rect 33 -1513 125 -1507
rect 191 -1473 283 -1467
rect 191 -1507 203 -1473
rect 271 -1507 283 -1473
rect 191 -1513 283 -1507
rect 349 -1473 441 -1467
rect 349 -1507 361 -1473
rect 429 -1507 441 -1473
rect 349 -1513 441 -1507
rect 507 -1473 599 -1467
rect 507 -1507 519 -1473
rect 587 -1507 599 -1473
rect 507 -1513 599 -1507
rect 665 -1473 757 -1467
rect 665 -1507 677 -1473
rect 745 -1507 757 -1473
rect 665 -1513 757 -1507
rect 823 -1473 915 -1467
rect 823 -1507 835 -1473
rect 903 -1507 915 -1473
rect 823 -1513 915 -1507
rect 981 -1473 1073 -1467
rect 981 -1507 993 -1473
rect 1061 -1507 1073 -1473
rect 981 -1513 1073 -1507
rect -1129 -1566 -1083 -1554
rect -1129 -2742 -1123 -1566
rect -1089 -2742 -1083 -1566
rect -1129 -2754 -1083 -2742
rect -971 -1566 -925 -1554
rect -971 -2742 -965 -1566
rect -931 -2742 -925 -1566
rect -971 -2754 -925 -2742
rect -813 -1566 -767 -1554
rect -813 -2742 -807 -1566
rect -773 -2742 -767 -1566
rect -813 -2754 -767 -2742
rect -655 -1566 -609 -1554
rect -655 -2742 -649 -1566
rect -615 -2742 -609 -1566
rect -655 -2754 -609 -2742
rect -497 -1566 -451 -1554
rect -497 -2742 -491 -1566
rect -457 -2742 -451 -1566
rect -497 -2754 -451 -2742
rect -339 -1566 -293 -1554
rect -339 -2742 -333 -1566
rect -299 -2742 -293 -1566
rect -339 -2754 -293 -2742
rect -181 -1566 -135 -1554
rect -181 -2742 -175 -1566
rect -141 -2742 -135 -1566
rect -181 -2754 -135 -2742
rect -23 -1566 23 -1554
rect -23 -2742 -17 -1566
rect 17 -2742 23 -1566
rect -23 -2754 23 -2742
rect 135 -1566 181 -1554
rect 135 -2742 141 -1566
rect 175 -2742 181 -1566
rect 135 -2754 181 -2742
rect 293 -1566 339 -1554
rect 293 -2742 299 -1566
rect 333 -2742 339 -1566
rect 293 -2754 339 -2742
rect 451 -1566 497 -1554
rect 451 -2742 457 -1566
rect 491 -2742 497 -1566
rect 451 -2754 497 -2742
rect 609 -1566 655 -1554
rect 609 -2742 615 -1566
rect 649 -2742 655 -1566
rect 609 -2754 655 -2742
rect 767 -1566 813 -1554
rect 767 -2742 773 -1566
rect 807 -2742 813 -1566
rect 767 -2754 813 -2742
rect 925 -1566 971 -1554
rect 925 -2742 931 -1566
rect 965 -2742 971 -1566
rect 925 -2754 971 -2742
rect 1083 -1566 1129 -1554
rect 1083 -2742 1089 -1566
rect 1123 -2742 1129 -1566
rect 1083 -2754 1129 -2742
rect -1073 -2801 -981 -2795
rect -1073 -2835 -1061 -2801
rect -993 -2835 -981 -2801
rect -1073 -2841 -981 -2835
rect -915 -2801 -823 -2795
rect -915 -2835 -903 -2801
rect -835 -2835 -823 -2801
rect -915 -2841 -823 -2835
rect -757 -2801 -665 -2795
rect -757 -2835 -745 -2801
rect -677 -2835 -665 -2801
rect -757 -2841 -665 -2835
rect -599 -2801 -507 -2795
rect -599 -2835 -587 -2801
rect -519 -2835 -507 -2801
rect -599 -2841 -507 -2835
rect -441 -2801 -349 -2795
rect -441 -2835 -429 -2801
rect -361 -2835 -349 -2801
rect -441 -2841 -349 -2835
rect -283 -2801 -191 -2795
rect -283 -2835 -271 -2801
rect -203 -2835 -191 -2801
rect -283 -2841 -191 -2835
rect -125 -2801 -33 -2795
rect -125 -2835 -113 -2801
rect -45 -2835 -33 -2801
rect -125 -2841 -33 -2835
rect 33 -2801 125 -2795
rect 33 -2835 45 -2801
rect 113 -2835 125 -2801
rect 33 -2841 125 -2835
rect 191 -2801 283 -2795
rect 191 -2835 203 -2801
rect 271 -2835 283 -2801
rect 191 -2841 283 -2835
rect 349 -2801 441 -2795
rect 349 -2835 361 -2801
rect 429 -2835 441 -2801
rect 349 -2841 441 -2835
rect 507 -2801 599 -2795
rect 507 -2835 519 -2801
rect 587 -2835 599 -2801
rect 507 -2841 599 -2835
rect 665 -2801 757 -2795
rect 665 -2835 677 -2801
rect 745 -2835 757 -2801
rect 665 -2841 757 -2835
rect 823 -2801 915 -2795
rect 823 -2835 835 -2801
rect 903 -2835 915 -2801
rect 823 -2841 915 -2835
rect 981 -2801 1073 -2795
rect 981 -2835 993 -2801
rect 1061 -2835 1073 -2801
rect 981 -2841 1073 -2835
<< properties >>
string FIXED_BBOX -1220 -2920 1220 2920
string gencell sky130_fd_pr__pfet_01v8_lvt
string library sky130
string parameters w 6.0 l 0.5 m 4 nf 14 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.35 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
