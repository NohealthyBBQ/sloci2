magic
tech sky130A
magscale 1 2
timestamp 1672344136
<< nwell >>
rect -1747 -984 1747 984
<< pmoslvt >>
rect -1551 -764 -1451 836
rect -1393 -764 -1293 836
rect -1235 -764 -1135 836
rect -1077 -764 -977 836
rect -919 -764 -819 836
rect -761 -764 -661 836
rect -603 -764 -503 836
rect -445 -764 -345 836
rect -287 -764 -187 836
rect -129 -764 -29 836
rect 29 -764 129 836
rect 187 -764 287 836
rect 345 -764 445 836
rect 503 -764 603 836
rect 661 -764 761 836
rect 819 -764 919 836
rect 977 -764 1077 836
rect 1135 -764 1235 836
rect 1293 -764 1393 836
rect 1451 -764 1551 836
<< pdiff >>
rect -1609 824 -1551 836
rect -1609 -752 -1597 824
rect -1563 -752 -1551 824
rect -1609 -764 -1551 -752
rect -1451 824 -1393 836
rect -1451 -752 -1439 824
rect -1405 -752 -1393 824
rect -1451 -764 -1393 -752
rect -1293 824 -1235 836
rect -1293 -752 -1281 824
rect -1247 -752 -1235 824
rect -1293 -764 -1235 -752
rect -1135 824 -1077 836
rect -1135 -752 -1123 824
rect -1089 -752 -1077 824
rect -1135 -764 -1077 -752
rect -977 824 -919 836
rect -977 -752 -965 824
rect -931 -752 -919 824
rect -977 -764 -919 -752
rect -819 824 -761 836
rect -819 -752 -807 824
rect -773 -752 -761 824
rect -819 -764 -761 -752
rect -661 824 -603 836
rect -661 -752 -649 824
rect -615 -752 -603 824
rect -661 -764 -603 -752
rect -503 824 -445 836
rect -503 -752 -491 824
rect -457 -752 -445 824
rect -503 -764 -445 -752
rect -345 824 -287 836
rect -345 -752 -333 824
rect -299 -752 -287 824
rect -345 -764 -287 -752
rect -187 824 -129 836
rect -187 -752 -175 824
rect -141 -752 -129 824
rect -187 -764 -129 -752
rect -29 824 29 836
rect -29 -752 -17 824
rect 17 -752 29 824
rect -29 -764 29 -752
rect 129 824 187 836
rect 129 -752 141 824
rect 175 -752 187 824
rect 129 -764 187 -752
rect 287 824 345 836
rect 287 -752 299 824
rect 333 -752 345 824
rect 287 -764 345 -752
rect 445 824 503 836
rect 445 -752 457 824
rect 491 -752 503 824
rect 445 -764 503 -752
rect 603 824 661 836
rect 603 -752 615 824
rect 649 -752 661 824
rect 603 -764 661 -752
rect 761 824 819 836
rect 761 -752 773 824
rect 807 -752 819 824
rect 761 -764 819 -752
rect 919 824 977 836
rect 919 -752 931 824
rect 965 -752 977 824
rect 919 -764 977 -752
rect 1077 824 1135 836
rect 1077 -752 1089 824
rect 1123 -752 1135 824
rect 1077 -764 1135 -752
rect 1235 824 1293 836
rect 1235 -752 1247 824
rect 1281 -752 1293 824
rect 1235 -764 1293 -752
rect 1393 824 1451 836
rect 1393 -752 1405 824
rect 1439 -752 1451 824
rect 1393 -764 1451 -752
rect 1551 824 1609 836
rect 1551 -752 1563 824
rect 1597 -752 1609 824
rect 1551 -764 1609 -752
<< pdiffc >>
rect -1597 -752 -1563 824
rect -1439 -752 -1405 824
rect -1281 -752 -1247 824
rect -1123 -752 -1089 824
rect -965 -752 -931 824
rect -807 -752 -773 824
rect -649 -752 -615 824
rect -491 -752 -457 824
rect -333 -752 -299 824
rect -175 -752 -141 824
rect -17 -752 17 824
rect 141 -752 175 824
rect 299 -752 333 824
rect 457 -752 491 824
rect 615 -752 649 824
rect 773 -752 807 824
rect 931 -752 965 824
rect 1089 -752 1123 824
rect 1247 -752 1281 824
rect 1405 -752 1439 824
rect 1563 -752 1597 824
<< nsubdiff >>
rect -1711 914 -1615 948
rect 1615 914 1711 948
rect -1711 851 -1677 914
rect 1677 851 1711 914
rect -1711 -914 -1677 -851
rect 1677 -914 1711 -851
rect -1711 -948 -1615 -914
rect 1615 -948 1711 -914
<< nsubdiffcont >>
rect -1615 914 1615 948
rect -1711 -851 -1677 851
rect 1677 -851 1711 851
rect -1615 -948 1615 -914
<< poly >>
rect -1551 836 -1451 862
rect -1393 836 -1293 862
rect -1235 836 -1135 862
rect -1077 836 -977 862
rect -919 836 -819 862
rect -761 836 -661 862
rect -603 836 -503 862
rect -445 836 -345 862
rect -287 836 -187 862
rect -129 836 -29 862
rect 29 836 129 862
rect 187 836 287 862
rect 345 836 445 862
rect 503 836 603 862
rect 661 836 761 862
rect 819 836 919 862
rect 977 836 1077 862
rect 1135 836 1235 862
rect 1293 836 1393 862
rect 1451 836 1551 862
rect -1551 -811 -1451 -764
rect -1551 -845 -1535 -811
rect -1467 -845 -1451 -811
rect -1551 -861 -1451 -845
rect -1393 -811 -1293 -764
rect -1393 -845 -1377 -811
rect -1309 -845 -1293 -811
rect -1393 -861 -1293 -845
rect -1235 -811 -1135 -764
rect -1235 -845 -1219 -811
rect -1151 -845 -1135 -811
rect -1235 -861 -1135 -845
rect -1077 -811 -977 -764
rect -1077 -845 -1061 -811
rect -993 -845 -977 -811
rect -1077 -861 -977 -845
rect -919 -811 -819 -764
rect -919 -845 -903 -811
rect -835 -845 -819 -811
rect -919 -861 -819 -845
rect -761 -811 -661 -764
rect -761 -845 -745 -811
rect -677 -845 -661 -811
rect -761 -861 -661 -845
rect -603 -811 -503 -764
rect -603 -845 -587 -811
rect -519 -845 -503 -811
rect -603 -861 -503 -845
rect -445 -811 -345 -764
rect -445 -845 -429 -811
rect -361 -845 -345 -811
rect -445 -861 -345 -845
rect -287 -811 -187 -764
rect -287 -845 -271 -811
rect -203 -845 -187 -811
rect -287 -861 -187 -845
rect -129 -811 -29 -764
rect -129 -845 -113 -811
rect -45 -845 -29 -811
rect -129 -861 -29 -845
rect 29 -811 129 -764
rect 29 -845 45 -811
rect 113 -845 129 -811
rect 29 -861 129 -845
rect 187 -811 287 -764
rect 187 -845 203 -811
rect 271 -845 287 -811
rect 187 -861 287 -845
rect 345 -811 445 -764
rect 345 -845 361 -811
rect 429 -845 445 -811
rect 345 -861 445 -845
rect 503 -811 603 -764
rect 503 -845 519 -811
rect 587 -845 603 -811
rect 503 -861 603 -845
rect 661 -811 761 -764
rect 661 -845 677 -811
rect 745 -845 761 -811
rect 661 -861 761 -845
rect 819 -811 919 -764
rect 819 -845 835 -811
rect 903 -845 919 -811
rect 819 -861 919 -845
rect 977 -811 1077 -764
rect 977 -845 993 -811
rect 1061 -845 1077 -811
rect 977 -861 1077 -845
rect 1135 -811 1235 -764
rect 1135 -845 1151 -811
rect 1219 -845 1235 -811
rect 1135 -861 1235 -845
rect 1293 -811 1393 -764
rect 1293 -845 1309 -811
rect 1377 -845 1393 -811
rect 1293 -861 1393 -845
rect 1451 -811 1551 -764
rect 1451 -845 1467 -811
rect 1535 -845 1551 -811
rect 1451 -861 1551 -845
<< polycont >>
rect -1535 -845 -1467 -811
rect -1377 -845 -1309 -811
rect -1219 -845 -1151 -811
rect -1061 -845 -993 -811
rect -903 -845 -835 -811
rect -745 -845 -677 -811
rect -587 -845 -519 -811
rect -429 -845 -361 -811
rect -271 -845 -203 -811
rect -113 -845 -45 -811
rect 45 -845 113 -811
rect 203 -845 271 -811
rect 361 -845 429 -811
rect 519 -845 587 -811
rect 677 -845 745 -811
rect 835 -845 903 -811
rect 993 -845 1061 -811
rect 1151 -845 1219 -811
rect 1309 -845 1377 -811
rect 1467 -845 1535 -811
<< locali >>
rect -1711 914 -1615 948
rect 1615 914 1711 948
rect -1711 851 -1677 914
rect 1677 851 1711 914
rect -1597 824 -1563 840
rect -1597 -768 -1563 -752
rect -1439 824 -1405 840
rect -1439 -768 -1405 -752
rect -1281 824 -1247 840
rect -1281 -768 -1247 -752
rect -1123 824 -1089 840
rect -1123 -768 -1089 -752
rect -965 824 -931 840
rect -965 -768 -931 -752
rect -807 824 -773 840
rect -807 -768 -773 -752
rect -649 824 -615 840
rect -649 -768 -615 -752
rect -491 824 -457 840
rect -491 -768 -457 -752
rect -333 824 -299 840
rect -333 -768 -299 -752
rect -175 824 -141 840
rect -175 -768 -141 -752
rect -17 824 17 840
rect -17 -768 17 -752
rect 141 824 175 840
rect 141 -768 175 -752
rect 299 824 333 840
rect 299 -768 333 -752
rect 457 824 491 840
rect 457 -768 491 -752
rect 615 824 649 840
rect 615 -768 649 -752
rect 773 824 807 840
rect 773 -768 807 -752
rect 931 824 965 840
rect 931 -768 965 -752
rect 1089 824 1123 840
rect 1089 -768 1123 -752
rect 1247 824 1281 840
rect 1247 -768 1281 -752
rect 1405 824 1439 840
rect 1405 -768 1439 -752
rect 1563 824 1597 840
rect 1563 -768 1597 -752
rect -1551 -845 -1535 -811
rect -1467 -845 -1451 -811
rect -1393 -845 -1377 -811
rect -1309 -845 -1293 -811
rect -1235 -845 -1219 -811
rect -1151 -845 -1135 -811
rect -1077 -845 -1061 -811
rect -993 -845 -977 -811
rect -919 -845 -903 -811
rect -835 -845 -819 -811
rect -761 -845 -745 -811
rect -677 -845 -661 -811
rect -603 -845 -587 -811
rect -519 -845 -503 -811
rect -445 -845 -429 -811
rect -361 -845 -345 -811
rect -287 -845 -271 -811
rect -203 -845 -187 -811
rect -129 -845 -113 -811
rect -45 -845 -29 -811
rect 29 -845 45 -811
rect 113 -845 129 -811
rect 187 -845 203 -811
rect 271 -845 287 -811
rect 345 -845 361 -811
rect 429 -845 445 -811
rect 503 -845 519 -811
rect 587 -845 603 -811
rect 661 -845 677 -811
rect 745 -845 761 -811
rect 819 -845 835 -811
rect 903 -845 919 -811
rect 977 -845 993 -811
rect 1061 -845 1077 -811
rect 1135 -845 1151 -811
rect 1219 -845 1235 -811
rect 1293 -845 1309 -811
rect 1377 -845 1393 -811
rect 1451 -845 1467 -811
rect 1535 -845 1551 -811
rect -1711 -914 -1677 -851
rect 1677 -914 1711 -851
rect -1711 -948 -1615 -914
rect 1615 -948 1711 -914
<< viali >>
rect -1597 -752 -1563 824
rect -1439 -752 -1405 824
rect -1281 -752 -1247 824
rect -1123 -752 -1089 824
rect -965 -752 -931 824
rect -807 -752 -773 824
rect -649 -752 -615 824
rect -491 -752 -457 824
rect -333 -752 -299 824
rect -175 -752 -141 824
rect -17 -752 17 824
rect 141 -752 175 824
rect 299 -752 333 824
rect 457 -752 491 824
rect 615 -752 649 824
rect 773 -752 807 824
rect 931 -752 965 824
rect 1089 -752 1123 824
rect 1247 -752 1281 824
rect 1405 -752 1439 824
rect 1563 -752 1597 824
rect -1535 -845 -1467 -811
rect -1377 -845 -1309 -811
rect -1219 -845 -1151 -811
rect -1061 -845 -993 -811
rect -903 -845 -835 -811
rect -745 -845 -677 -811
rect -587 -845 -519 -811
rect -429 -845 -361 -811
rect -271 -845 -203 -811
rect -113 -845 -45 -811
rect 45 -845 113 -811
rect 203 -845 271 -811
rect 361 -845 429 -811
rect 519 -845 587 -811
rect 677 -845 745 -811
rect 835 -845 903 -811
rect 993 -845 1061 -811
rect 1151 -845 1219 -811
rect 1309 -845 1377 -811
rect 1467 -845 1535 -811
<< metal1 >>
rect -1603 824 -1557 836
rect -1603 -752 -1597 824
rect -1563 -752 -1557 824
rect -1603 -764 -1557 -752
rect -1445 824 -1399 836
rect -1445 -752 -1439 824
rect -1405 -752 -1399 824
rect -1445 -764 -1399 -752
rect -1287 824 -1241 836
rect -1287 -752 -1281 824
rect -1247 -752 -1241 824
rect -1287 -764 -1241 -752
rect -1129 824 -1083 836
rect -1129 -752 -1123 824
rect -1089 -752 -1083 824
rect -1129 -764 -1083 -752
rect -971 824 -925 836
rect -971 -752 -965 824
rect -931 -752 -925 824
rect -971 -764 -925 -752
rect -813 824 -767 836
rect -813 -752 -807 824
rect -773 -752 -767 824
rect -813 -764 -767 -752
rect -655 824 -609 836
rect -655 -752 -649 824
rect -615 -752 -609 824
rect -655 -764 -609 -752
rect -497 824 -451 836
rect -497 -752 -491 824
rect -457 -752 -451 824
rect -497 -764 -451 -752
rect -339 824 -293 836
rect -339 -752 -333 824
rect -299 -752 -293 824
rect -339 -764 -293 -752
rect -181 824 -135 836
rect -181 -752 -175 824
rect -141 -752 -135 824
rect -181 -764 -135 -752
rect -23 824 23 836
rect -23 -752 -17 824
rect 17 -752 23 824
rect -23 -764 23 -752
rect 135 824 181 836
rect 135 -752 141 824
rect 175 -752 181 824
rect 135 -764 181 -752
rect 293 824 339 836
rect 293 -752 299 824
rect 333 -752 339 824
rect 293 -764 339 -752
rect 451 824 497 836
rect 451 -752 457 824
rect 491 -752 497 824
rect 451 -764 497 -752
rect 609 824 655 836
rect 609 -752 615 824
rect 649 -752 655 824
rect 609 -764 655 -752
rect 767 824 813 836
rect 767 -752 773 824
rect 807 -752 813 824
rect 767 -764 813 -752
rect 925 824 971 836
rect 925 -752 931 824
rect 965 -752 971 824
rect 925 -764 971 -752
rect 1083 824 1129 836
rect 1083 -752 1089 824
rect 1123 -752 1129 824
rect 1083 -764 1129 -752
rect 1241 824 1287 836
rect 1241 -752 1247 824
rect 1281 -752 1287 824
rect 1241 -764 1287 -752
rect 1399 824 1445 836
rect 1399 -752 1405 824
rect 1439 -752 1445 824
rect 1399 -764 1445 -752
rect 1557 824 1603 836
rect 1557 -752 1563 824
rect 1597 -752 1603 824
rect 1557 -764 1603 -752
rect -1547 -811 -1455 -805
rect -1547 -845 -1535 -811
rect -1467 -845 -1455 -811
rect -1547 -851 -1455 -845
rect -1389 -811 -1297 -805
rect -1389 -845 -1377 -811
rect -1309 -845 -1297 -811
rect -1389 -851 -1297 -845
rect -1231 -811 -1139 -805
rect -1231 -845 -1219 -811
rect -1151 -845 -1139 -811
rect -1231 -851 -1139 -845
rect -1073 -811 -981 -805
rect -1073 -845 -1061 -811
rect -993 -845 -981 -811
rect -1073 -851 -981 -845
rect -915 -811 -823 -805
rect -915 -845 -903 -811
rect -835 -845 -823 -811
rect -915 -851 -823 -845
rect -757 -811 -665 -805
rect -757 -845 -745 -811
rect -677 -845 -665 -811
rect -757 -851 -665 -845
rect -599 -811 -507 -805
rect -599 -845 -587 -811
rect -519 -845 -507 -811
rect -599 -851 -507 -845
rect -441 -811 -349 -805
rect -441 -845 -429 -811
rect -361 -845 -349 -811
rect -441 -851 -349 -845
rect -283 -811 -191 -805
rect -283 -845 -271 -811
rect -203 -845 -191 -811
rect -283 -851 -191 -845
rect -125 -811 -33 -805
rect -125 -845 -113 -811
rect -45 -845 -33 -811
rect -125 -851 -33 -845
rect 33 -811 125 -805
rect 33 -845 45 -811
rect 113 -845 125 -811
rect 33 -851 125 -845
rect 191 -811 283 -805
rect 191 -845 203 -811
rect 271 -845 283 -811
rect 191 -851 283 -845
rect 349 -811 441 -805
rect 349 -845 361 -811
rect 429 -845 441 -811
rect 349 -851 441 -845
rect 507 -811 599 -805
rect 507 -845 519 -811
rect 587 -845 599 -811
rect 507 -851 599 -845
rect 665 -811 757 -805
rect 665 -845 677 -811
rect 745 -845 757 -811
rect 665 -851 757 -845
rect 823 -811 915 -805
rect 823 -845 835 -811
rect 903 -845 915 -811
rect 823 -851 915 -845
rect 981 -811 1073 -805
rect 981 -845 993 -811
rect 1061 -845 1073 -811
rect 981 -851 1073 -845
rect 1139 -811 1231 -805
rect 1139 -845 1151 -811
rect 1219 -845 1231 -811
rect 1139 -851 1231 -845
rect 1297 -811 1389 -805
rect 1297 -845 1309 -811
rect 1377 -845 1389 -811
rect 1297 -851 1389 -845
rect 1455 -811 1547 -805
rect 1455 -845 1467 -811
rect 1535 -845 1547 -811
rect 1455 -851 1547 -845
<< properties >>
string FIXED_BBOX -1694 -931 1694 931
string gencell sky130_fd_pr__pfet_01v8_lvt
string library sky130
string parameters w 8 l 0.5 m 1 nf 20 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 0 botc 1 poverlap 0 doverlap 1 lmin 0.35 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
