magic
tech sky130A
magscale 1 2
timestamp 1662515374
<< pwell >>
rect 4320 3755 4385 3760
rect 2396 3114 2534 3552
rect 4195 1515 4300 1600
rect 4405 1400 4510 1410
rect 4205 1315 4295 1400
rect 4180 1120 4190 1210
<< locali >>
rect 3915 3945 4040 3980
rect 3265 3645 3380 3680
rect 4580 3650 4730 3685
rect 3260 3335 3385 3370
rect 3920 3335 4045 3370
rect 4580 3335 4705 3370
rect 3260 3185 3385 3220
rect 3890 3185 4070 3220
rect 4550 3185 4705 3220
rect 2435 2260 2470 2460
rect 3265 1035 3390 1070
rect 3920 1035 4045 1070
rect 4580 1035 4705 1070
<< metal1 >>
rect 3550 3890 3635 3900
rect 3550 3820 3560 3890
rect 3625 3820 3635 3890
rect 4325 3890 4410 3900
rect 3640 3868 3750 3874
rect 3738 3834 3750 3868
rect 3640 3828 3750 3834
rect 3780 3835 3875 3845
rect 3550 3810 3635 3820
rect 3665 3790 3750 3800
rect 3665 3778 3675 3790
rect 3550 3772 3675 3778
rect 3425 3735 3520 3745
rect 3425 3675 3435 3735
rect 3490 3675 3520 3735
rect 3550 3738 3562 3772
rect 3665 3738 3675 3772
rect 3550 3732 3675 3738
rect 3665 3720 3675 3732
rect 3740 3720 3750 3790
rect 3780 3775 3810 3835
rect 3865 3775 3875 3835
rect 3780 3765 3875 3775
rect 4085 3835 4180 3845
rect 4085 3775 4095 3835
rect 4150 3775 4180 3835
rect 4325 3820 4335 3890
rect 4400 3820 4410 3890
rect 4325 3810 4410 3820
rect 4085 3765 4180 3775
rect 4210 3790 4295 3800
rect 3665 3710 3750 3720
rect 4210 3720 4220 3790
rect 4285 3720 4295 3790
rect 4210 3710 4295 3720
rect 4440 3735 4535 3745
rect 3425 3665 3520 3675
rect 3550 3690 3635 3700
rect 3550 3625 3560 3690
rect 3625 3682 3635 3690
rect 4325 3690 4410 3700
rect 3625 3676 3750 3682
rect 3625 3642 3635 3676
rect 3738 3642 3750 3676
rect 3625 3636 3750 3642
rect 3780 3640 3875 3650
rect 3625 3625 3635 3636
rect 3550 3615 3635 3625
rect 3665 3595 3750 3605
rect 3665 3586 3675 3595
rect 3550 3580 3675 3586
rect 3425 3545 3520 3555
rect 3425 3485 3435 3545
rect 3490 3485 3520 3545
rect 3550 3546 3562 3580
rect 3665 3546 3675 3580
rect 3550 3540 3675 3546
rect 3665 3530 3675 3540
rect 3740 3530 3750 3595
rect 3780 3580 3810 3640
rect 3865 3580 3875 3640
rect 3780 3570 3875 3580
rect 4085 3640 4180 3650
rect 4085 3580 4095 3640
rect 4150 3580 4180 3640
rect 4325 3625 4335 3690
rect 4400 3625 4410 3690
rect 4440 3675 4470 3735
rect 4525 3675 4535 3735
rect 4440 3665 4535 3675
rect 4325 3615 4410 3625
rect 4085 3570 4180 3580
rect 4210 3595 4295 3605
rect 3665 3520 3750 3530
rect 4210 3530 4220 3595
rect 4285 3530 4295 3595
rect 4210 3520 4295 3530
rect 4440 3545 4535 3555
rect 3425 3475 3520 3485
rect 3550 3500 3635 3510
rect 3550 3430 3560 3500
rect 3625 3490 3635 3500
rect 4325 3500 4410 3510
rect 3625 3484 3750 3490
rect 3625 3450 3635 3484
rect 3738 3450 3750 3484
rect 3625 3444 3750 3450
rect 3625 3430 3635 3444
rect 3550 3420 3635 3430
rect 4325 3430 4335 3500
rect 4400 3430 4410 3500
rect 4440 3485 4470 3545
rect 4525 3485 4535 3545
rect 4440 3475 4535 3485
rect 4325 3420 4410 3430
rect 3665 3125 3750 3135
rect 3665 3110 3675 3125
rect 3550 3103 3675 3110
rect 3550 3070 3562 3103
rect 3665 3070 3675 3103
rect 3550 3063 3675 3070
rect 3665 3060 3675 3063
rect 3740 3060 3750 3125
rect 4210 3125 4295 3135
rect 3665 3050 3750 3060
rect 3780 3070 3875 3080
rect 3550 3025 3635 3035
rect 3425 2970 3520 2980
rect 3425 2910 3435 2970
rect 3490 2910 3520 2970
rect 3550 2960 3560 3025
rect 3625 3014 3635 3025
rect 3625 3007 3750 3014
rect 3625 2974 3635 3007
rect 3738 2974 3750 3007
rect 3780 3010 3810 3070
rect 3865 3010 3875 3070
rect 3780 3000 3875 3010
rect 4085 3070 4180 3080
rect 4085 3010 4095 3070
rect 4150 3010 4180 3070
rect 4210 3060 4220 3125
rect 4285 3110 4295 3125
rect 4285 3103 4410 3110
rect 4285 3070 4295 3103
rect 4398 3070 4410 3103
rect 4285 3063 4410 3070
rect 4285 3060 4295 3063
rect 4210 3050 4295 3060
rect 4325 3025 4410 3035
rect 4325 3014 4335 3025
rect 4085 3000 4180 3010
rect 4210 3007 4335 3014
rect 3625 2967 3750 2974
rect 4210 2974 4222 3007
rect 4325 2974 4335 3007
rect 4210 2967 4335 2974
rect 3625 2960 3635 2967
rect 3550 2950 3635 2960
rect 4325 2960 4335 2967
rect 4400 2960 4410 3025
rect 4325 2950 4410 2960
rect 4440 2970 4535 2980
rect 3665 2925 3750 2935
rect 3665 2918 3675 2925
rect 3425 2900 3520 2910
rect 3550 2911 3675 2918
rect 3550 2878 3562 2911
rect 3665 2878 3675 2911
rect 3550 2871 3675 2878
rect 3665 2860 3675 2871
rect 3740 2860 3750 2925
rect 4210 2925 4295 2935
rect 3665 2850 3750 2860
rect 3780 2875 3875 2885
rect 3550 2830 3635 2840
rect 3425 2780 3520 2790
rect 3425 2720 3435 2780
rect 3490 2720 3520 2780
rect 3550 2765 3560 2830
rect 3625 2822 3635 2830
rect 3625 2815 3750 2822
rect 3625 2782 3635 2815
rect 3738 2782 3750 2815
rect 3780 2815 3810 2875
rect 3865 2815 3875 2875
rect 3780 2805 3875 2815
rect 4085 2875 4180 2885
rect 4085 2815 4095 2875
rect 4150 2815 4180 2875
rect 4210 2860 4220 2925
rect 4285 2918 4295 2925
rect 4285 2911 4410 2918
rect 4285 2878 4295 2911
rect 4398 2878 4410 2911
rect 4440 2910 4470 2970
rect 4525 2910 4535 2970
rect 4440 2900 4535 2910
rect 4285 2871 4410 2878
rect 4285 2860 4295 2871
rect 4210 2850 4295 2860
rect 4325 2830 4410 2840
rect 4325 2822 4335 2830
rect 4085 2805 4180 2815
rect 4210 2815 4335 2822
rect 3625 2775 3750 2782
rect 4210 2782 4222 2815
rect 4325 2782 4335 2815
rect 4210 2775 4335 2782
rect 3625 2765 3635 2775
rect 3550 2755 3635 2765
rect 4325 2765 4335 2775
rect 4400 2765 4410 2830
rect 4325 2755 4410 2765
rect 4440 2780 4535 2790
rect 3665 2735 3750 2745
rect 3665 2726 3675 2735
rect 3425 2710 3520 2720
rect 3550 2718 3675 2726
rect 3550 2686 3562 2718
rect 3665 2686 3675 2718
rect 3550 2678 3675 2686
rect 3665 2675 3675 2678
rect 3740 2675 3750 2735
rect 4210 2735 4295 2745
rect 3665 2665 3750 2675
rect 3780 2685 3875 2695
rect 3550 2640 3635 2650
rect 3425 2590 3520 2600
rect 3425 2530 3435 2590
rect 3490 2530 3520 2590
rect 3550 2575 3560 2640
rect 3625 2630 3635 2640
rect 3625 2622 3750 2630
rect 3625 2590 3635 2622
rect 3738 2590 3750 2622
rect 3780 2625 3810 2685
rect 3865 2625 3875 2685
rect 3780 2615 3875 2625
rect 4085 2685 4180 2695
rect 4085 2625 4095 2685
rect 4150 2625 4180 2685
rect 4210 2675 4220 2735
rect 4285 2726 4295 2735
rect 4285 2718 4410 2726
rect 4285 2686 4295 2718
rect 4398 2686 4410 2718
rect 4440 2720 4470 2780
rect 4525 2720 4535 2780
rect 4440 2710 4535 2720
rect 4285 2678 4410 2686
rect 4285 2675 4295 2678
rect 4210 2665 4295 2675
rect 4325 2640 4410 2650
rect 4325 2630 4335 2640
rect 4085 2615 4180 2625
rect 4210 2622 4335 2630
rect 3625 2582 3750 2590
rect 4210 2590 4222 2622
rect 4325 2590 4335 2622
rect 4210 2582 4335 2590
rect 3625 2575 3635 2582
rect 3550 2565 3635 2575
rect 4325 2575 4335 2582
rect 4400 2575 4410 2640
rect 4325 2565 4410 2575
rect 4440 2590 4535 2600
rect 3665 2540 3750 2550
rect 3665 2534 3675 2540
rect 3425 2520 3520 2530
rect 3550 2526 3675 2534
rect 3550 2494 3562 2526
rect 3665 2494 3675 2526
rect 3550 2486 3675 2494
rect 3665 2480 3675 2486
rect 3740 2480 3750 2540
rect 4210 2540 4295 2550
rect 3665 2470 3750 2480
rect 3780 2490 3875 2500
rect 3550 2445 3635 2455
rect 3425 2400 3520 2410
rect 3425 2340 3435 2400
rect 3490 2340 3520 2400
rect 3550 2385 3560 2445
rect 3625 2438 3635 2445
rect 3625 2430 3750 2438
rect 3625 2398 3635 2430
rect 3738 2398 3750 2430
rect 3780 2430 3810 2490
rect 3865 2430 3875 2490
rect 3780 2420 3875 2430
rect 4085 2490 4180 2500
rect 4085 2430 4095 2490
rect 4150 2430 4180 2490
rect 4210 2480 4220 2540
rect 4285 2534 4295 2540
rect 4285 2526 4410 2534
rect 4285 2494 4295 2526
rect 4398 2494 4410 2526
rect 4440 2530 4470 2590
rect 4525 2530 4535 2590
rect 4440 2520 4535 2530
rect 4285 2486 4410 2494
rect 4285 2480 4295 2486
rect 4210 2470 4295 2480
rect 4325 2445 4410 2455
rect 4325 2438 4335 2445
rect 4085 2420 4180 2430
rect 4210 2430 4335 2438
rect 3625 2390 3750 2398
rect 4210 2398 4222 2430
rect 4325 2398 4335 2430
rect 4210 2390 4335 2398
rect 3625 2385 3635 2390
rect 3550 2375 3635 2385
rect 4325 2385 4335 2390
rect 4400 2385 4410 2445
rect 4325 2375 4410 2385
rect 4440 2400 4535 2410
rect 3665 2350 3750 2360
rect 3665 2344 3675 2350
rect 3425 2330 3520 2340
rect 3550 2336 3675 2344
rect 3550 2304 3562 2336
rect 3665 2304 3675 2336
rect 3550 2296 3675 2304
rect 3665 2290 3675 2296
rect 3740 2290 3750 2350
rect 4210 2350 4295 2360
rect 3665 2280 3750 2290
rect 3780 2300 3875 2310
rect 3550 2255 3635 2265
rect 3425 2205 3520 2215
rect 3425 2145 3435 2205
rect 3490 2145 3520 2205
rect 3550 2190 3560 2255
rect 3625 2248 3635 2255
rect 3625 2240 3750 2248
rect 3625 2208 3635 2240
rect 3738 2208 3750 2240
rect 3780 2240 3810 2300
rect 3865 2240 3875 2300
rect 3780 2230 3875 2240
rect 4085 2300 4180 2310
rect 4085 2240 4095 2300
rect 4150 2240 4180 2300
rect 4210 2290 4220 2350
rect 4285 2344 4295 2350
rect 4285 2336 4410 2344
rect 4285 2304 4295 2336
rect 4398 2304 4410 2336
rect 4440 2340 4470 2400
rect 4525 2340 4535 2400
rect 4440 2330 4535 2340
rect 4285 2296 4410 2304
rect 4285 2290 4295 2296
rect 4210 2280 4295 2290
rect 4325 2255 4410 2265
rect 4325 2248 4335 2255
rect 4085 2230 4180 2240
rect 4210 2240 4335 2248
rect 3625 2200 3750 2208
rect 4210 2208 4222 2240
rect 4325 2208 4335 2240
rect 4210 2200 4335 2208
rect 3625 2190 3635 2200
rect 3550 2180 3635 2190
rect 4325 2190 4335 2200
rect 4400 2190 4410 2255
rect 4325 2180 4410 2190
rect 4440 2205 4535 2215
rect 3665 2160 3750 2170
rect 3665 2152 3675 2160
rect 3425 2135 3520 2145
rect 3550 2144 3675 2152
rect 3550 2112 3562 2144
rect 3665 2112 3675 2144
rect 3550 2104 3675 2112
rect 3665 2095 3675 2104
rect 3740 2095 3750 2160
rect 4210 2160 4295 2170
rect 3665 2085 3750 2095
rect 3780 2110 3875 2120
rect 3550 2065 3635 2075
rect 3425 2015 3520 2025
rect 3425 1955 3435 2015
rect 3490 1955 3520 2015
rect 3550 2000 3560 2065
rect 3625 2056 3635 2065
rect 3625 2048 3750 2056
rect 3625 2016 3635 2048
rect 3738 2016 3750 2048
rect 3780 2050 3810 2110
rect 3865 2050 3875 2110
rect 3780 2040 3875 2050
rect 4085 2110 4180 2120
rect 4085 2050 4095 2110
rect 4150 2050 4180 2110
rect 4210 2095 4220 2160
rect 4285 2152 4295 2160
rect 4285 2144 4410 2152
rect 4285 2112 4295 2144
rect 4398 2112 4410 2144
rect 4440 2145 4470 2205
rect 4525 2145 4535 2205
rect 4440 2135 4535 2145
rect 4285 2104 4410 2112
rect 4285 2095 4295 2104
rect 4210 2085 4295 2095
rect 4325 2065 4410 2075
rect 4325 2056 4335 2065
rect 4085 2040 4180 2050
rect 4210 2048 4335 2056
rect 3625 2008 3750 2016
rect 4210 2016 4222 2048
rect 4325 2016 4335 2048
rect 4210 2008 4335 2016
rect 3625 2000 3635 2008
rect 3550 1990 3635 2000
rect 4325 2000 4335 2008
rect 4400 2000 4410 2065
rect 4325 1990 4410 2000
rect 4440 2015 4535 2025
rect 3665 1970 3750 1980
rect 3665 1959 3675 1970
rect 3425 1945 3520 1955
rect 3550 1952 3675 1959
rect 3550 1919 3562 1952
rect 3665 1919 3675 1952
rect 3550 1912 3675 1919
rect 3665 1905 3675 1912
rect 3740 1905 3750 1970
rect 4210 1970 4295 1980
rect 3665 1895 3750 1905
rect 3780 1915 3875 1925
rect 3550 1870 3635 1880
rect 3425 1820 3520 1830
rect 3425 1760 3435 1820
rect 3490 1760 3520 1820
rect 3550 1805 3560 1870
rect 3625 1863 3635 1870
rect 3625 1856 3750 1863
rect 3625 1823 3635 1856
rect 3738 1823 3750 1856
rect 3780 1855 3810 1915
rect 3865 1855 3875 1915
rect 3780 1845 3875 1855
rect 4085 1915 4180 1925
rect 4085 1855 4095 1915
rect 4150 1855 4180 1915
rect 4210 1905 4220 1970
rect 4285 1959 4295 1970
rect 4285 1952 4410 1959
rect 4285 1919 4295 1952
rect 4398 1919 4410 1952
rect 4440 1955 4470 2015
rect 4525 1955 4535 2015
rect 4440 1945 4535 1955
rect 4285 1912 4410 1919
rect 4285 1905 4295 1912
rect 4210 1895 4295 1905
rect 4325 1870 4410 1880
rect 4325 1863 4335 1870
rect 4085 1845 4180 1855
rect 4210 1856 4335 1863
rect 3625 1816 3750 1823
rect 4210 1823 4222 1856
rect 4325 1823 4335 1856
rect 4210 1816 4335 1823
rect 3625 1805 3635 1816
rect 3550 1795 3635 1805
rect 4325 1805 4335 1816
rect 4400 1805 4410 1870
rect 4325 1795 4410 1805
rect 4440 1820 4535 1830
rect 3665 1775 3750 1785
rect 3665 1767 3675 1775
rect 3425 1750 3520 1760
rect 3550 1760 3675 1767
rect 3550 1727 3562 1760
rect 3665 1727 3675 1760
rect 3550 1720 3675 1727
rect 3665 1710 3675 1720
rect 3740 1710 3750 1775
rect 4210 1775 4295 1785
rect 3665 1700 3750 1710
rect 3780 1725 3875 1735
rect 3550 1680 3635 1690
rect 3425 1630 3520 1640
rect 2565 1580 3135 1600
rect 2565 1185 2585 1580
rect 3115 1185 3135 1580
rect 3425 1570 3435 1630
rect 3490 1570 3520 1630
rect 3550 1615 3560 1680
rect 3625 1671 3635 1680
rect 3625 1664 3750 1671
rect 3625 1631 3635 1664
rect 3738 1631 3750 1664
rect 3780 1665 3810 1725
rect 3865 1665 3875 1725
rect 3780 1655 3875 1665
rect 4085 1725 4180 1735
rect 4085 1665 4095 1725
rect 4150 1665 4180 1725
rect 4210 1710 4220 1775
rect 4285 1767 4295 1775
rect 4285 1760 4410 1767
rect 4285 1727 4295 1760
rect 4398 1727 4410 1760
rect 4440 1760 4470 1820
rect 4525 1760 4535 1820
rect 4440 1750 4535 1760
rect 4285 1720 4410 1727
rect 4285 1710 4295 1720
rect 4210 1700 4295 1710
rect 4325 1680 4410 1690
rect 4325 1671 4335 1680
rect 4085 1655 4180 1665
rect 4210 1664 4335 1671
rect 3625 1624 3750 1631
rect 4210 1631 4222 1664
rect 4325 1631 4335 1664
rect 4210 1624 4335 1631
rect 3625 1615 3635 1624
rect 3550 1605 3635 1615
rect 4325 1615 4335 1624
rect 4400 1615 4410 1680
rect 4325 1605 4410 1615
rect 4440 1630 4535 1640
rect 3665 1585 3750 1595
rect 3665 1574 3675 1585
rect 3425 1560 3520 1570
rect 3550 1568 3675 1574
rect 3550 1534 3562 1568
rect 3665 1534 3675 1568
rect 3550 1528 3675 1534
rect 3665 1520 3675 1528
rect 3740 1520 3750 1585
rect 4210 1585 4295 1595
rect 3665 1510 3750 1520
rect 3780 1530 3875 1540
rect 3550 1485 3635 1500
rect 3425 1435 3520 1445
rect 3425 1375 3435 1435
rect 3490 1375 3520 1435
rect 3550 1420 3560 1485
rect 3625 1478 3635 1485
rect 3625 1472 3750 1478
rect 3625 1438 3635 1472
rect 3738 1438 3750 1472
rect 3780 1470 3810 1530
rect 3865 1470 3875 1530
rect 3780 1460 3875 1470
rect 4085 1530 4180 1540
rect 4085 1470 4095 1530
rect 4150 1470 4180 1530
rect 4210 1520 4220 1585
rect 4285 1574 4295 1585
rect 4285 1568 4410 1574
rect 4285 1534 4295 1568
rect 4398 1534 4410 1568
rect 4440 1570 4470 1630
rect 4525 1570 4535 1630
rect 4440 1560 4535 1570
rect 4825 1580 5395 1600
rect 4285 1528 4410 1534
rect 4285 1520 4295 1528
rect 4210 1510 4295 1520
rect 4325 1485 4410 1500
rect 4325 1478 4335 1485
rect 4085 1460 4180 1470
rect 4210 1472 4335 1478
rect 3625 1432 3750 1438
rect 4210 1438 4222 1472
rect 4325 1438 4335 1472
rect 4210 1432 4335 1438
rect 3625 1420 3635 1432
rect 3550 1410 3635 1420
rect 4325 1420 4335 1432
rect 4400 1420 4410 1485
rect 4325 1410 4410 1420
rect 4440 1435 4535 1445
rect 3665 1390 3750 1400
rect 3665 1382 3675 1390
rect 3425 1365 3520 1375
rect 3550 1376 3675 1382
rect 3550 1342 3562 1376
rect 3665 1342 3675 1376
rect 3550 1336 3675 1342
rect 3665 1325 3675 1336
rect 3740 1325 3750 1390
rect 4210 1390 4295 1400
rect 3665 1315 3750 1325
rect 3780 1340 3875 1350
rect 3550 1295 3635 1305
rect 2565 1165 3135 1185
rect 3425 1245 3520 1255
rect 3425 1185 3435 1245
rect 3490 1185 3520 1245
rect 3550 1230 3560 1295
rect 3625 1286 3635 1295
rect 3625 1280 3750 1286
rect 3625 1246 3635 1280
rect 3738 1246 3750 1280
rect 3780 1280 3810 1340
rect 3865 1280 3875 1340
rect 3780 1270 3875 1280
rect 4085 1340 4180 1350
rect 4085 1280 4095 1340
rect 4150 1280 4180 1340
rect 4210 1325 4220 1390
rect 4285 1382 4295 1390
rect 4285 1376 4410 1382
rect 4285 1342 4295 1376
rect 4398 1342 4410 1376
rect 4440 1375 4470 1435
rect 4525 1375 4535 1435
rect 4440 1365 4535 1375
rect 4285 1336 4410 1342
rect 4285 1325 4295 1336
rect 4210 1315 4295 1325
rect 4325 1295 4410 1305
rect 4325 1286 4335 1295
rect 4085 1270 4180 1280
rect 4210 1280 4335 1286
rect 3625 1240 3750 1246
rect 4210 1246 4222 1280
rect 4325 1246 4335 1280
rect 4210 1240 4335 1246
rect 3625 1230 3635 1240
rect 3550 1220 3635 1230
rect 4325 1230 4335 1240
rect 4400 1230 4410 1295
rect 4325 1220 4410 1230
rect 4440 1245 4535 1255
rect 3665 1200 3750 1210
rect 3665 1190 3675 1200
rect 3425 1175 3520 1185
rect 3550 1184 3675 1190
rect 3550 1150 3562 1184
rect 3665 1150 3675 1184
rect 3550 1144 3675 1150
rect 3665 1130 3675 1144
rect 3740 1130 3750 1200
rect 3665 1120 3750 1130
rect 4210 1200 4295 1210
rect 4210 1130 4220 1200
rect 4285 1190 4295 1200
rect 4285 1184 4410 1190
rect 4285 1150 4295 1184
rect 4398 1150 4410 1184
rect 4440 1185 4470 1245
rect 4525 1185 4535 1245
rect 4440 1175 4535 1185
rect 4825 1185 4845 1580
rect 5375 1185 5395 1580
rect 4825 1165 5395 1185
rect 4285 1144 4410 1150
rect 4285 1130 4295 1144
rect 4210 1120 4295 1130
<< via1 >>
rect 3560 3820 3625 3890
rect 3435 3675 3490 3735
rect 3675 3720 3740 3790
rect 3810 3775 3865 3835
rect 4095 3775 4150 3835
rect 4335 3820 4400 3890
rect 4220 3720 4285 3790
rect 3560 3625 3625 3690
rect 2585 3140 3115 3530
rect 3435 3485 3490 3545
rect 3675 3530 3740 3595
rect 3810 3580 3865 3640
rect 4095 3580 4150 3640
rect 4335 3625 4400 3690
rect 4470 3675 4525 3735
rect 4220 3530 4285 3595
rect 3560 3430 3625 3500
rect 4335 3430 4400 3500
rect 4470 3485 4525 3545
rect 4845 3140 5375 3530
rect 3675 3060 3740 3125
rect 3435 2910 3490 2970
rect 3560 2960 3625 3025
rect 3810 3010 3865 3070
rect 4095 3010 4150 3070
rect 4220 3060 4285 3125
rect 4335 2960 4400 3025
rect 3675 2860 3740 2925
rect 3435 2720 3490 2780
rect 3560 2765 3625 2830
rect 3810 2815 3865 2875
rect 4095 2815 4150 2875
rect 4220 2860 4285 2925
rect 4470 2910 4525 2970
rect 4335 2765 4400 2830
rect 3675 2675 3740 2735
rect 3435 2530 3490 2590
rect 3560 2575 3625 2640
rect 3810 2625 3865 2685
rect 4095 2625 4150 2685
rect 4220 2675 4285 2735
rect 4470 2720 4525 2780
rect 4335 2575 4400 2640
rect 3675 2480 3740 2540
rect 3435 2340 3490 2400
rect 3560 2385 3625 2445
rect 3810 2430 3865 2490
rect 4095 2430 4150 2490
rect 4220 2480 4285 2540
rect 4470 2530 4525 2590
rect 4335 2385 4400 2445
rect 3675 2290 3740 2350
rect 3435 2145 3490 2205
rect 3560 2190 3625 2255
rect 3810 2240 3865 2300
rect 4095 2240 4150 2300
rect 4220 2290 4285 2350
rect 4470 2340 4525 2400
rect 4335 2190 4400 2255
rect 3675 2095 3740 2160
rect 3435 1955 3490 2015
rect 3560 2000 3625 2065
rect 3810 2050 3865 2110
rect 4095 2050 4150 2110
rect 4220 2095 4285 2160
rect 4470 2145 4525 2205
rect 4335 2000 4400 2065
rect 3675 1905 3740 1970
rect 3435 1760 3490 1820
rect 3560 1805 3625 1870
rect 3810 1855 3865 1915
rect 4095 1855 4150 1915
rect 4220 1905 4285 1970
rect 4470 1955 4525 2015
rect 4335 1805 4400 1870
rect 3675 1710 3740 1775
rect 2585 1185 3115 1580
rect 3435 1570 3490 1630
rect 3560 1615 3625 1680
rect 3810 1665 3865 1725
rect 4095 1665 4150 1725
rect 4220 1710 4285 1775
rect 4470 1760 4525 1820
rect 4335 1615 4400 1680
rect 3675 1520 3740 1585
rect 3435 1375 3490 1435
rect 3560 1420 3625 1485
rect 3810 1470 3865 1530
rect 4095 1470 4150 1530
rect 4220 1520 4285 1585
rect 4470 1570 4525 1630
rect 4335 1420 4400 1485
rect 3675 1325 3740 1390
rect 3435 1185 3490 1245
rect 3560 1230 3625 1295
rect 3810 1280 3865 1340
rect 4095 1280 4150 1340
rect 4220 1325 4285 1390
rect 4470 1375 4525 1435
rect 4335 1230 4400 1295
rect 3675 1130 3740 1200
rect 4220 1130 4285 1200
rect 4470 1185 4525 1245
rect 4845 1185 5375 1580
<< metal2 >>
rect 3425 3945 3875 4020
rect 3425 3735 3500 3945
rect 3530 3890 3635 3900
rect 3530 3820 3540 3890
rect 3625 3820 3635 3890
rect 3530 3810 3635 3820
rect 3800 3835 3875 3945
rect 3425 3675 3435 3735
rect 3490 3675 3500 3735
rect 3665 3790 3770 3800
rect 3665 3720 3675 3790
rect 3760 3720 3770 3790
rect 3665 3710 3770 3720
rect 3800 3775 3810 3835
rect 3865 3775 3875 3835
rect 2565 3530 3135 3550
rect 2565 3140 2585 3530
rect 3115 3140 3135 3530
rect 3425 3545 3500 3675
rect 3530 3690 3635 3700
rect 3530 3625 3540 3690
rect 3625 3625 3635 3690
rect 3530 3615 3635 3625
rect 3800 3640 3875 3775
rect 3425 3485 3435 3545
rect 3490 3485 3500 3545
rect 3665 3595 3770 3605
rect 3665 3530 3675 3595
rect 3760 3530 3770 3595
rect 3800 3580 3810 3640
rect 3865 3580 3875 3640
rect 3800 3570 3875 3580
rect 4085 3945 4535 4020
rect 4085 3835 4160 3945
rect 4085 3775 4095 3835
rect 4150 3775 4160 3835
rect 4325 3890 4430 3900
rect 4325 3820 4335 3890
rect 4420 3820 4430 3890
rect 4325 3810 4430 3820
rect 4085 3640 4160 3775
rect 4190 3790 4295 3800
rect 4190 3720 4200 3790
rect 4285 3720 4295 3790
rect 4190 3710 4295 3720
rect 4460 3735 4535 3945
rect 4085 3580 4095 3640
rect 4150 3580 4160 3640
rect 4325 3690 4430 3700
rect 4325 3625 4335 3690
rect 4420 3625 4430 3690
rect 4325 3615 4430 3625
rect 4460 3675 4470 3735
rect 4525 3675 4535 3735
rect 4085 3570 4160 3580
rect 4190 3595 4295 3605
rect 3665 3520 3770 3530
rect 4190 3530 4200 3595
rect 4285 3530 4295 3595
rect 4190 3520 4295 3530
rect 4460 3545 4535 3675
rect 3425 3475 3500 3485
rect 3530 3500 3635 3510
rect 3530 3430 3540 3500
rect 3625 3430 3635 3500
rect 3530 3420 3635 3430
rect 4325 3500 4430 3510
rect 4325 3430 4335 3500
rect 4420 3430 4430 3500
rect 4460 3485 4470 3545
rect 4525 3485 4535 3545
rect 4460 3475 4535 3485
rect 4825 3530 5395 3550
rect 4325 3420 4430 3430
rect 2565 3120 3135 3140
rect 4825 3140 4845 3530
rect 5375 3140 5395 3530
rect 3665 3125 3770 3135
rect 3665 3060 3675 3125
rect 3760 3060 3770 3125
rect 4190 3125 4295 3135
rect 3665 3050 3770 3060
rect 3800 3070 3875 3080
rect 3535 3025 3635 3035
rect 3425 2970 3500 2980
rect 3425 2910 3435 2970
rect 3490 2910 3500 2970
rect 3535 2960 3540 3025
rect 3625 2960 3635 3025
rect 3535 2950 3635 2960
rect 3800 3010 3810 3070
rect 3865 3010 3875 3070
rect 3425 2780 3500 2910
rect 3665 2925 3770 2935
rect 3665 2860 3675 2925
rect 3760 2860 3770 2925
rect 3665 2850 3770 2860
rect 3800 2875 3875 3010
rect 3425 2720 3435 2780
rect 3490 2720 3500 2780
rect 3535 2830 3635 2840
rect 3535 2765 3540 2830
rect 3625 2765 3635 2830
rect 3535 2755 3635 2765
rect 3800 2815 3810 2875
rect 3865 2815 3875 2875
rect 3425 2590 3500 2720
rect 3665 2735 3770 2750
rect 3665 2675 3675 2735
rect 3760 2675 3770 2735
rect 3665 2665 3770 2675
rect 3800 2685 3875 2815
rect 3425 2530 3435 2590
rect 3490 2530 3500 2590
rect 3535 2640 3635 2650
rect 3535 2575 3540 2640
rect 3625 2575 3635 2640
rect 3535 2565 3635 2575
rect 3800 2625 3810 2685
rect 3865 2625 3875 2685
rect 3425 2400 3500 2530
rect 3665 2540 3770 2550
rect 3665 2480 3675 2540
rect 3760 2480 3770 2540
rect 3665 2470 3770 2480
rect 3800 2490 3875 2625
rect 3425 2340 3435 2400
rect 3490 2340 3500 2400
rect 3535 2445 3635 2455
rect 3535 2385 3540 2445
rect 3625 2385 3635 2445
rect 3535 2375 3635 2385
rect 3800 2430 3810 2490
rect 3865 2430 3875 2490
rect 3425 2205 3500 2340
rect 3665 2350 3770 2365
rect 3665 2290 3675 2350
rect 3760 2290 3770 2350
rect 3665 2280 3770 2290
rect 3800 2300 3875 2430
rect 3425 2145 3435 2205
rect 3490 2145 3500 2205
rect 3535 2255 3635 2265
rect 3535 2190 3540 2255
rect 3625 2190 3635 2255
rect 3535 2180 3635 2190
rect 3800 2240 3810 2300
rect 3865 2240 3875 2300
rect 3425 2015 3500 2145
rect 3665 2160 3770 2170
rect 3665 2095 3675 2160
rect 3760 2095 3770 2160
rect 3665 2085 3770 2095
rect 3800 2110 3875 2240
rect 3425 1955 3435 2015
rect 3490 1955 3500 2015
rect 3535 2065 3635 2075
rect 3535 2000 3540 2065
rect 3625 2000 3635 2065
rect 3535 1990 3635 2000
rect 3800 2050 3810 2110
rect 3865 2050 3875 2110
rect 3425 1820 3500 1955
rect 3665 1970 3770 1980
rect 3665 1905 3675 1970
rect 3760 1905 3770 1970
rect 3665 1895 3770 1905
rect 3800 1915 3875 2050
rect 3425 1760 3435 1820
rect 3490 1760 3500 1820
rect 3535 1870 3635 1880
rect 3535 1805 3540 1870
rect 3625 1805 3635 1870
rect 3535 1795 3635 1805
rect 3800 1855 3810 1915
rect 3865 1855 3875 1915
rect 3425 1630 3500 1760
rect 3665 1775 3770 1785
rect 3665 1710 3675 1775
rect 3760 1710 3770 1775
rect 3665 1700 3770 1710
rect 3800 1725 3875 1855
rect 2565 1580 3135 1600
rect 2565 1185 2585 1580
rect 3115 1185 3135 1580
rect 2565 610 3135 1185
rect 2565 355 2585 610
rect 3115 355 3135 610
rect 2565 335 3135 355
rect 3425 1570 3435 1630
rect 3490 1570 3500 1630
rect 3535 1680 3635 1690
rect 3535 1615 3540 1680
rect 3625 1615 3635 1680
rect 3535 1605 3635 1615
rect 3800 1665 3810 1725
rect 3865 1665 3875 1725
rect 3425 1435 3500 1570
rect 3665 1585 3770 1595
rect 3665 1520 3675 1585
rect 3760 1520 3770 1585
rect 3665 1510 3770 1520
rect 3800 1530 3875 1665
rect 3425 1375 3435 1435
rect 3490 1375 3500 1435
rect 3535 1485 3635 1495
rect 3535 1420 3540 1485
rect 3625 1420 3635 1485
rect 3535 1410 3635 1420
rect 3800 1470 3810 1530
rect 3865 1470 3875 1530
rect 3425 1245 3500 1375
rect 3665 1390 3770 1400
rect 3665 1325 3675 1390
rect 3760 1325 3770 1390
rect 3665 1315 3770 1325
rect 3800 1340 3875 1470
rect 3425 1185 3435 1245
rect 3490 1185 3500 1245
rect 3530 1295 3635 1305
rect 3530 1230 3540 1295
rect 3625 1230 3635 1295
rect 3530 1220 3635 1230
rect 3800 1280 3810 1340
rect 3865 1280 3875 1340
rect 3425 305 3500 1185
rect 3665 1200 3770 1210
rect 3665 1130 3675 1200
rect 3760 1130 3770 1200
rect 3665 1120 3770 1130
rect 3800 305 3875 1280
rect 4085 3070 4160 3080
rect 4085 3010 4095 3070
rect 4150 3010 4160 3070
rect 4190 3060 4200 3125
rect 4285 3060 4295 3125
rect 4825 3120 5395 3140
rect 4190 3050 4295 3060
rect 4085 2875 4160 3010
rect 4325 3025 4425 3035
rect 4325 2960 4335 3025
rect 4420 2960 4425 3025
rect 4325 2950 4425 2960
rect 4460 2970 4535 2980
rect 4085 2815 4095 2875
rect 4150 2815 4160 2875
rect 4190 2925 4295 2935
rect 4190 2860 4200 2925
rect 4285 2860 4295 2925
rect 4190 2850 4295 2860
rect 4460 2910 4470 2970
rect 4525 2910 4535 2970
rect 4085 2685 4160 2815
rect 4325 2830 4425 2840
rect 4325 2765 4335 2830
rect 4420 2765 4425 2830
rect 4325 2755 4425 2765
rect 4460 2780 4535 2910
rect 4085 2625 4095 2685
rect 4150 2625 4160 2685
rect 4190 2735 4295 2750
rect 4190 2675 4200 2735
rect 4285 2675 4295 2735
rect 4190 2665 4295 2675
rect 4460 2720 4470 2780
rect 4525 2720 4535 2780
rect 4085 2490 4160 2625
rect 4325 2640 4425 2650
rect 4325 2575 4335 2640
rect 4420 2575 4425 2640
rect 4325 2565 4425 2575
rect 4460 2590 4535 2720
rect 4085 2430 4095 2490
rect 4150 2430 4160 2490
rect 4190 2540 4295 2550
rect 4190 2480 4200 2540
rect 4285 2480 4295 2540
rect 4190 2470 4295 2480
rect 4460 2530 4470 2590
rect 4525 2530 4535 2590
rect 4085 2300 4160 2430
rect 4325 2445 4425 2455
rect 4325 2385 4335 2445
rect 4420 2385 4425 2445
rect 4325 2375 4425 2385
rect 4460 2400 4535 2530
rect 4085 2240 4095 2300
rect 4150 2240 4160 2300
rect 4190 2350 4295 2365
rect 4190 2290 4200 2350
rect 4285 2290 4295 2350
rect 4190 2280 4295 2290
rect 4460 2340 4470 2400
rect 4525 2340 4535 2400
rect 4085 2110 4160 2240
rect 4325 2255 4425 2265
rect 4325 2190 4335 2255
rect 4420 2190 4425 2255
rect 4325 2180 4425 2190
rect 4460 2205 4535 2340
rect 4085 2050 4095 2110
rect 4150 2050 4160 2110
rect 4190 2160 4295 2170
rect 4190 2095 4200 2160
rect 4285 2095 4295 2160
rect 4190 2085 4295 2095
rect 4460 2145 4470 2205
rect 4525 2145 4535 2205
rect 4085 1915 4160 2050
rect 4325 2065 4425 2075
rect 4325 2000 4335 2065
rect 4420 2000 4425 2065
rect 4325 1990 4425 2000
rect 4460 2015 4535 2145
rect 4085 1855 4095 1915
rect 4150 1855 4160 1915
rect 4190 1970 4295 1980
rect 4190 1905 4200 1970
rect 4285 1905 4295 1970
rect 4190 1895 4295 1905
rect 4460 1955 4470 2015
rect 4525 1955 4535 2015
rect 4085 1725 4160 1855
rect 4325 1870 4425 1880
rect 4325 1805 4335 1870
rect 4420 1805 4425 1870
rect 4325 1795 4425 1805
rect 4460 1820 4535 1955
rect 4085 1665 4095 1725
rect 4150 1665 4160 1725
rect 4190 1775 4295 1785
rect 4190 1710 4200 1775
rect 4285 1710 4295 1775
rect 4190 1700 4295 1710
rect 4460 1760 4470 1820
rect 4525 1760 4535 1820
rect 4085 1530 4160 1665
rect 4325 1680 4425 1690
rect 4325 1615 4335 1680
rect 4420 1615 4425 1680
rect 4325 1605 4425 1615
rect 4460 1630 4535 1760
rect 4085 1470 4095 1530
rect 4150 1470 4160 1530
rect 4190 1585 4295 1595
rect 4190 1520 4200 1585
rect 4285 1520 4295 1585
rect 4190 1510 4295 1520
rect 4460 1570 4470 1630
rect 4525 1570 4535 1630
rect 4085 1340 4160 1470
rect 4325 1485 4425 1495
rect 4325 1420 4335 1485
rect 4420 1420 4425 1485
rect 4325 1410 4425 1420
rect 4460 1435 4535 1570
rect 4085 1280 4095 1340
rect 4150 1280 4160 1340
rect 4190 1390 4295 1400
rect 4190 1325 4200 1390
rect 4285 1325 4295 1390
rect 4190 1315 4295 1325
rect 4460 1375 4470 1435
rect 4525 1375 4535 1435
rect 4085 305 4160 1280
rect 4325 1295 4430 1305
rect 4325 1230 4335 1295
rect 4420 1230 4430 1295
rect 4325 1220 4430 1230
rect 4460 1245 4535 1375
rect 4190 1200 4295 1210
rect 4190 1130 4200 1200
rect 4285 1130 4295 1200
rect 4190 1120 4295 1130
rect 4460 1185 4470 1245
rect 4525 1185 4535 1245
rect 4460 305 4535 1185
rect 4825 1580 5395 1600
rect 4825 1185 4845 1580
rect 5375 1185 5395 1580
rect 4825 615 5395 1185
rect 4825 355 4845 615
rect 5375 355 5395 615
rect 4825 335 5395 355
rect 2400 230 4535 305
<< via2 >>
rect 3540 3820 3560 3890
rect 3560 3820 3610 3890
rect 3690 3720 3740 3790
rect 3740 3720 3760 3790
rect 2585 3140 3115 3530
rect 3540 3625 3560 3690
rect 3560 3625 3610 3690
rect 3690 3530 3740 3595
rect 3740 3530 3760 3595
rect 4350 3820 4400 3890
rect 4400 3820 4420 3890
rect 4200 3720 4220 3790
rect 4220 3720 4270 3790
rect 4350 3625 4400 3690
rect 4400 3625 4420 3690
rect 4200 3530 4220 3595
rect 4220 3530 4270 3595
rect 3540 3430 3560 3500
rect 3560 3430 3610 3500
rect 4350 3430 4400 3500
rect 4400 3430 4420 3500
rect 4845 3140 5375 3530
rect 3690 3060 3740 3125
rect 3740 3060 3760 3125
rect 3540 2960 3560 3025
rect 3560 2960 3610 3025
rect 3690 2860 3740 2925
rect 3740 2860 3760 2925
rect 3540 2765 3560 2830
rect 3560 2765 3610 2830
rect 3690 2675 3740 2735
rect 3740 2675 3760 2735
rect 3540 2575 3560 2640
rect 3560 2575 3610 2640
rect 3690 2480 3740 2540
rect 3740 2480 3760 2540
rect 3540 2385 3560 2445
rect 3560 2385 3610 2445
rect 3690 2290 3740 2350
rect 3740 2290 3760 2350
rect 3540 2190 3560 2255
rect 3560 2190 3610 2255
rect 3690 2095 3740 2160
rect 3740 2095 3760 2160
rect 3540 2000 3560 2065
rect 3560 2000 3610 2065
rect 3690 1905 3740 1970
rect 3740 1905 3760 1970
rect 3540 1805 3560 1870
rect 3560 1805 3610 1870
rect 3690 1710 3740 1775
rect 3740 1710 3760 1775
rect 2585 355 3115 610
rect 3540 1615 3560 1680
rect 3560 1615 3610 1680
rect 3690 1520 3740 1585
rect 3740 1520 3760 1585
rect 3540 1420 3560 1485
rect 3560 1420 3610 1485
rect 3690 1325 3740 1390
rect 3740 1325 3760 1390
rect 3540 1230 3560 1295
rect 3560 1230 3610 1295
rect 3690 1130 3740 1200
rect 3740 1130 3760 1200
rect 4200 3060 4220 3125
rect 4220 3060 4270 3125
rect 4350 2960 4400 3025
rect 4400 2960 4420 3025
rect 4200 2860 4220 2925
rect 4220 2860 4270 2925
rect 4350 2765 4400 2830
rect 4400 2765 4420 2830
rect 4200 2675 4220 2735
rect 4220 2675 4270 2735
rect 4350 2575 4400 2640
rect 4400 2575 4420 2640
rect 4200 2480 4220 2540
rect 4220 2480 4270 2540
rect 4350 2385 4400 2445
rect 4400 2385 4420 2445
rect 4200 2290 4220 2350
rect 4220 2290 4270 2350
rect 4350 2190 4400 2255
rect 4400 2190 4420 2255
rect 4200 2095 4220 2160
rect 4220 2095 4270 2160
rect 4350 2000 4400 2065
rect 4400 2000 4420 2065
rect 4200 1905 4220 1970
rect 4220 1905 4270 1970
rect 4350 1805 4400 1870
rect 4400 1805 4420 1870
rect 4200 1710 4220 1775
rect 4220 1710 4270 1775
rect 4350 1615 4400 1680
rect 4400 1615 4420 1680
rect 4200 1520 4220 1585
rect 4220 1520 4270 1585
rect 4350 1420 4400 1485
rect 4400 1420 4420 1485
rect 4200 1325 4220 1390
rect 4220 1325 4270 1390
rect 4350 1230 4400 1295
rect 4400 1230 4420 1295
rect 4200 1130 4220 1200
rect 4220 1130 4270 1200
rect 4845 355 5375 615
<< metal3 >>
rect 3320 3890 3620 3900
rect 3320 3820 3540 3890
rect 3610 3820 3620 3890
rect 4340 3890 4640 3900
rect 3320 3690 3620 3820
rect 3320 3625 3540 3690
rect 3610 3625 3620 3690
rect 3320 3600 3620 3625
rect 2566 3530 3620 3600
rect 2566 3140 2585 3530
rect 3115 3500 3620 3530
rect 3115 3430 3540 3500
rect 3610 3430 3620 3500
rect 3115 3300 3620 3430
rect 3680 3790 4280 3845
rect 3680 3720 3690 3790
rect 3760 3720 4200 3790
rect 4270 3720 4280 3790
rect 3680 3595 4280 3720
rect 3680 3530 3690 3595
rect 3760 3530 4200 3595
rect 4270 3530 4280 3595
rect 3115 3140 3135 3300
rect 3680 3155 4280 3530
rect 4340 3820 4350 3890
rect 4420 3820 4640 3890
rect 4340 3690 4640 3820
rect 4340 3625 4350 3690
rect 4420 3625 4640 3690
rect 4340 3600 4640 3625
rect 4340 3550 5395 3600
rect 4340 3530 5396 3550
rect 4340 3500 4845 3530
rect 4340 3430 4350 3500
rect 4420 3430 4845 3500
rect 4340 3300 4845 3430
rect 2566 3120 3135 3140
rect 3320 3025 3620 3140
rect 3320 2960 3540 3025
rect 3610 2960 3620 3025
rect 3320 2830 3620 2960
rect 3320 2765 3540 2830
rect 3610 2765 3620 2830
rect 3320 2640 3620 2765
rect 3320 2575 3540 2640
rect 3610 2575 3620 2640
rect 3320 2445 3620 2575
rect 3320 2385 3540 2445
rect 3610 2385 3620 2445
rect 3320 2255 3620 2385
rect 3320 2190 3540 2255
rect 3610 2190 3620 2255
rect 3320 2065 3620 2190
rect 3320 2000 3540 2065
rect 3610 2000 3620 2065
rect 3320 1870 3620 2000
rect 3320 1805 3540 1870
rect 3610 1805 3620 1870
rect 3320 1680 3620 1805
rect 3320 1615 3540 1680
rect 3610 1615 3620 1680
rect 3320 1485 3620 1615
rect 3320 1420 3540 1485
rect 3610 1420 3620 1485
rect 3320 1295 3620 1420
rect 3320 1230 3540 1295
rect 3610 1230 3620 1295
rect 3320 1045 3620 1230
rect 3680 3125 3800 3155
rect 3680 3060 3690 3125
rect 3760 3080 3800 3125
rect 3875 3125 4280 3155
rect 4825 3140 4845 3300
rect 5375 3140 5396 3530
rect 3875 3080 4200 3125
rect 3760 3060 4200 3080
rect 4270 3060 4280 3125
rect 3680 2925 4280 3060
rect 3680 2860 3690 2925
rect 3760 2860 4200 2925
rect 4270 2860 4280 2925
rect 3680 2735 4280 2860
rect 3680 2675 3690 2735
rect 3760 2675 4200 2735
rect 4270 2675 4280 2735
rect 3680 2540 4280 2675
rect 3680 2480 3690 2540
rect 3760 2480 4200 2540
rect 4270 2480 4280 2540
rect 3680 2350 4280 2480
rect 3680 2290 3690 2350
rect 3760 2290 4200 2350
rect 4270 2290 4280 2350
rect 3680 2160 4280 2290
rect 3680 2095 3690 2160
rect 3760 2095 4200 2160
rect 4270 2095 4280 2160
rect 3680 1970 4280 2095
rect 3680 1905 3690 1970
rect 3760 1905 4200 1970
rect 4270 1905 4280 1970
rect 3680 1775 4280 1905
rect 3680 1710 3690 1775
rect 3760 1710 4200 1775
rect 4270 1710 4280 1775
rect 3680 1585 4280 1710
rect 3680 1520 3690 1585
rect 3760 1520 4200 1585
rect 4270 1520 4280 1585
rect 3680 1390 4280 1520
rect 3680 1325 3690 1390
rect 3760 1325 4200 1390
rect 4270 1325 4280 1390
rect 3680 1200 4280 1325
rect 3680 1130 3690 1200
rect 3760 1130 4200 1200
rect 4270 1130 4280 1200
rect 3680 1105 4280 1130
rect 4340 3025 4640 3140
rect 4825 3120 5396 3140
rect 4340 2960 4350 3025
rect 4420 2960 4640 3025
rect 4340 2830 4640 2960
rect 4340 2765 4350 2830
rect 4420 2765 4640 2830
rect 4340 2640 4640 2765
rect 4340 2575 4350 2640
rect 4420 2575 4640 2640
rect 4340 2445 4640 2575
rect 4340 2385 4350 2445
rect 4420 2385 4640 2445
rect 4340 2255 4640 2385
rect 4340 2190 4350 2255
rect 4420 2190 4640 2255
rect 4340 2065 4640 2190
rect 4340 2000 4350 2065
rect 4420 2000 4640 2065
rect 4340 1870 4640 2000
rect 4340 1805 4350 1870
rect 4420 1805 4640 1870
rect 4340 1680 4640 1805
rect 4340 1615 4350 1680
rect 4420 1615 4640 1680
rect 4340 1485 4640 1615
rect 4340 1420 4350 1485
rect 4420 1420 4640 1485
rect 4340 1295 4640 1420
rect 4340 1230 4350 1295
rect 4420 1230 4640 1295
rect 4340 1045 4640 1230
rect 2400 745 4640 1045
rect 2400 695 2700 745
rect 2400 615 5395 635
rect 2400 610 4845 615
rect 2400 355 2585 610
rect 3115 355 4845 610
rect 5375 355 5395 615
rect 2400 335 5395 355
use sky130_fd_pr__nfet_01v8_lvt_YTLFGX  XM1
timestamp 1662510845
transform 0 -1 3650 -1 0 2127
box -1127 -310 1127 310
use sky130_fd_pr__nfet_01v8_lvt_HNLS5R  XM2
timestamp 1662515274
transform 0 -1 3650 -1 0 3659
box -359 -310 359 310
use sky130_fd_pr__nfet_01v8_lvt_HNLS5R  XM3
timestamp 1662515274
transform 0 1 4310 -1 0 3659
box -359 -310 359 310
use sky130_fd_pr__nfet_01v8_lvt_YTLFGX  XM4
timestamp 1662510845
transform 0 1 4310 -1 0 2127
box -1127 -310 1127 310
use sky130_fd_pr__res_high_po_2p85_P79JE3  XR16
timestamp 1662404926
transform 1 0 2851 0 1 2358
box -451 -1358 451 1358
use sky130_fd_pr__res_high_po_2p85_P79JE3  XR17
timestamp 1662404926
transform 1 0 5111 0 1 2358
box -451 -1358 451 1358
<< labels >>
flabel metal2 3622 4000 3622 4000 1 FreeMono 2 0 0 0 INA
flabel metal2 4308 3992 4308 3992 1 FreeMono 2 0 0 0 INB
flabel metal3 2466 480 2466 480 1 FreeMono 2 0 0 0 VDD
flabel metal2 2472 260 2472 260 1 FreeMono 2 0 0 0 BIAS
rlabel metal2 2400 230 2514 304 1 BIAS
rlabel space 2398 336 2496 632 1 VDD
rlabel space 2396 700 2542 1048 1 GND
rlabel space 2430 2258 2468 2466 1 SUB
rlabel metal2 2400 230 4535 305 0 BIAS
rlabel metal3 2400 335 2585 635 0 VDD
rlabel metal3 2400 695 2700 1045 0 GND
rlabel metal2 3425 3945 3875 4020 1 INA
rlabel metal2 4085 3945 4535 4020 1 INB
rlabel locali 2435 2260 2470 2460 1 SUB
rlabel metal3 2566 3552 3136 3598 1 OUTA
rlabel metal3 4340 3530 5395 3600 1 OUTB
<< end >>
