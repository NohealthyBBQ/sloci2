magic
tech sky130A
magscale 1 2
timestamp 1662764279
<< nwell >>
rect -812 -284 812 284
<< pmoslvt >>
rect -616 -136 -416 64
rect -358 -136 -158 64
rect -100 -136 100 64
rect 158 -136 358 64
rect 416 -136 616 64
<< pdiff >>
rect -674 52 -616 64
rect -674 -124 -662 52
rect -628 -124 -616 52
rect -674 -136 -616 -124
rect -416 52 -358 64
rect -416 -124 -404 52
rect -370 -124 -358 52
rect -416 -136 -358 -124
rect -158 52 -100 64
rect -158 -124 -146 52
rect -112 -124 -100 52
rect -158 -136 -100 -124
rect 100 52 158 64
rect 100 -124 112 52
rect 146 -124 158 52
rect 100 -136 158 -124
rect 358 52 416 64
rect 358 -124 370 52
rect 404 -124 416 52
rect 358 -136 416 -124
rect 616 52 674 64
rect 616 -124 628 52
rect 662 -124 674 52
rect 616 -136 674 -124
<< pdiffc >>
rect -662 -124 -628 52
rect -404 -124 -370 52
rect -146 -124 -112 52
rect 112 -124 146 52
rect 370 -124 404 52
rect 628 -124 662 52
<< nsubdiff >>
rect -776 214 776 248
rect -776 151 -742 214
rect 742 151 776 214
rect -776 -214 -742 -151
rect 742 -214 776 -151
rect -776 -248 776 -214
<< nsubdiffcont >>
rect -776 -151 -742 151
rect 742 -151 776 151
<< poly >>
rect -616 145 -416 161
rect -616 111 -600 145
rect -432 111 -416 145
rect -616 64 -416 111
rect -358 145 -158 161
rect -358 111 -342 145
rect -174 111 -158 145
rect -358 64 -158 111
rect -100 145 100 161
rect -100 111 -84 145
rect 84 111 100 145
rect -100 64 100 111
rect 158 145 358 161
rect 158 111 174 145
rect 342 111 358 145
rect 158 64 358 111
rect 416 145 616 161
rect 416 111 432 145
rect 600 111 616 145
rect 416 64 616 111
rect -616 -162 -416 -136
rect -358 -162 -158 -136
rect -100 -162 100 -136
rect 158 -162 358 -136
rect 416 -162 616 -136
<< polycont >>
rect -600 111 -432 145
rect -342 111 -174 145
rect -84 111 84 145
rect 174 111 342 145
rect 432 111 600 145
<< locali >>
rect -776 214 776 248
rect -776 151 -742 214
rect 742 151 776 214
rect -616 111 -600 145
rect -432 111 -416 145
rect -358 111 -342 145
rect -174 111 -158 145
rect -100 111 -84 145
rect 84 111 100 145
rect 158 111 174 145
rect 342 111 358 145
rect 416 111 432 145
rect 600 111 616 145
rect -662 52 -628 68
rect -662 -140 -628 -124
rect -404 52 -370 68
rect -404 -140 -370 -124
rect -146 52 -112 68
rect -146 -140 -112 -124
rect 112 52 146 68
rect 112 -140 146 -124
rect 370 52 404 68
rect 370 -140 404 -124
rect 628 52 662 68
rect 628 -140 662 -124
rect -776 -214 -742 -151
rect 742 -214 776 -151
rect -776 -248 776 -214
<< viali >>
rect -600 111 -432 145
rect -342 111 -174 145
rect -84 111 84 145
rect 174 111 342 145
rect 432 111 600 145
rect -662 -124 -628 52
rect -404 -124 -370 52
rect -146 -124 -112 52
rect 112 -124 146 52
rect 370 -124 404 52
rect 628 -124 662 52
<< metal1 >>
rect -612 145 -420 151
rect -612 111 -600 145
rect -432 111 -420 145
rect -612 105 -420 111
rect -354 145 -162 151
rect -354 111 -342 145
rect -174 111 -162 145
rect -354 105 -162 111
rect -96 145 96 151
rect -96 111 -84 145
rect 84 111 96 145
rect -96 105 96 111
rect 162 145 354 151
rect 162 111 174 145
rect 342 111 354 145
rect 162 105 354 111
rect 420 145 612 151
rect 420 111 432 145
rect 600 111 612 145
rect 420 105 612 111
rect -668 52 -622 64
rect -668 -124 -662 52
rect -628 -124 -622 52
rect -668 -136 -622 -124
rect -410 52 -364 64
rect -410 -124 -404 52
rect -370 -124 -364 52
rect -410 -136 -364 -124
rect -152 52 -106 64
rect -152 -124 -146 52
rect -112 -124 -106 52
rect -152 -136 -106 -124
rect 106 52 152 64
rect 106 -124 112 52
rect 146 -124 152 52
rect 106 -136 152 -124
rect 364 52 410 64
rect 364 -124 370 52
rect 404 -124 410 52
rect 364 -136 410 -124
rect 622 52 668 64
rect 622 -124 628 52
rect 662 -124 668 52
rect 622 -136 668 -124
<< properties >>
string FIXED_BBOX -759 -231 759 231
string gencell sky130_fd_pr__pfet_01v8_lvt
string library sky130
string parameters w 1 l 1 m 1 nf 5 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 0 gbc 0 tbcov 100 rlcov 100 topc 1 botc 0 poverlap 0 doverlap 1 lmin 0.35 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
