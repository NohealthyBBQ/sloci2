magic
tech sky130A
magscale 1 2
timestamp 1672262880
<< pwell >>
rect -2686 -279 2686 279
<< nmoslvt >>
rect -2490 -131 -2090 69
rect -2032 -131 -1632 69
rect -1574 -131 -1174 69
rect -1116 -131 -716 69
rect -658 -131 -258 69
rect -200 -131 200 69
rect 258 -131 658 69
rect 716 -131 1116 69
rect 1174 -131 1574 69
rect 1632 -131 2032 69
rect 2090 -131 2490 69
<< ndiff >>
rect -2548 57 -2490 69
rect -2548 -119 -2536 57
rect -2502 -119 -2490 57
rect -2548 -131 -2490 -119
rect -2090 57 -2032 69
rect -2090 -119 -2078 57
rect -2044 -119 -2032 57
rect -2090 -131 -2032 -119
rect -1632 57 -1574 69
rect -1632 -119 -1620 57
rect -1586 -119 -1574 57
rect -1632 -131 -1574 -119
rect -1174 57 -1116 69
rect -1174 -119 -1162 57
rect -1128 -119 -1116 57
rect -1174 -131 -1116 -119
rect -716 57 -658 69
rect -716 -119 -704 57
rect -670 -119 -658 57
rect -716 -131 -658 -119
rect -258 57 -200 69
rect -258 -119 -246 57
rect -212 -119 -200 57
rect -258 -131 -200 -119
rect 200 57 258 69
rect 200 -119 212 57
rect 246 -119 258 57
rect 200 -131 258 -119
rect 658 57 716 69
rect 658 -119 670 57
rect 704 -119 716 57
rect 658 -131 716 -119
rect 1116 57 1174 69
rect 1116 -119 1128 57
rect 1162 -119 1174 57
rect 1116 -131 1174 -119
rect 1574 57 1632 69
rect 1574 -119 1586 57
rect 1620 -119 1632 57
rect 1574 -131 1632 -119
rect 2032 57 2090 69
rect 2032 -119 2044 57
rect 2078 -119 2090 57
rect 2032 -131 2090 -119
rect 2490 57 2548 69
rect 2490 -119 2502 57
rect 2536 -119 2548 57
rect 2490 -131 2548 -119
<< ndiffc >>
rect -2536 -119 -2502 57
rect -2078 -119 -2044 57
rect -1620 -119 -1586 57
rect -1162 -119 -1128 57
rect -704 -119 -670 57
rect -246 -119 -212 57
rect 212 -119 246 57
rect 670 -119 704 57
rect 1128 -119 1162 57
rect 1586 -119 1620 57
rect 2044 -119 2078 57
rect 2502 -119 2536 57
<< psubdiff >>
rect -2650 209 -2554 243
rect 2554 209 2650 243
rect -2650 -209 -2616 209
rect 2616 -209 2650 209
rect -2650 -243 2650 -209
<< psubdiffcont >>
rect -2554 209 2554 243
<< poly >>
rect -2490 141 -2090 157
rect -2490 107 -2474 141
rect -2106 107 -2090 141
rect -2490 69 -2090 107
rect -2032 141 -1632 157
rect -2032 107 -2016 141
rect -1648 107 -1632 141
rect -2032 69 -1632 107
rect -1574 141 -1174 157
rect -1574 107 -1558 141
rect -1190 107 -1174 141
rect -1574 69 -1174 107
rect -1116 141 -716 157
rect -1116 107 -1100 141
rect -732 107 -716 141
rect -1116 69 -716 107
rect -658 141 -258 157
rect -658 107 -642 141
rect -274 107 -258 141
rect -658 69 -258 107
rect -200 141 200 157
rect -200 107 -184 141
rect 184 107 200 141
rect -200 69 200 107
rect 258 141 658 157
rect 258 107 274 141
rect 642 107 658 141
rect 258 69 658 107
rect 716 141 1116 157
rect 716 107 732 141
rect 1100 107 1116 141
rect 716 69 1116 107
rect 1174 141 1574 157
rect 1174 107 1190 141
rect 1558 107 1574 141
rect 1174 69 1574 107
rect 1632 141 2032 157
rect 1632 107 1648 141
rect 2016 107 2032 141
rect 1632 69 2032 107
rect 2090 141 2490 157
rect 2090 107 2106 141
rect 2474 107 2490 141
rect 2090 69 2490 107
rect -2490 -157 -2090 -131
rect -2032 -157 -1632 -131
rect -1574 -157 -1174 -131
rect -1116 -157 -716 -131
rect -658 -157 -258 -131
rect -200 -157 200 -131
rect 258 -157 658 -131
rect 716 -157 1116 -131
rect 1174 -157 1574 -131
rect 1632 -157 2032 -131
rect 2090 -157 2490 -131
<< polycont >>
rect -2474 107 -2106 141
rect -2016 107 -1648 141
rect -1558 107 -1190 141
rect -1100 107 -732 141
rect -642 107 -274 141
rect -184 107 184 141
rect 274 107 642 141
rect 732 107 1100 141
rect 1190 107 1558 141
rect 1648 107 2016 141
rect 2106 107 2474 141
<< locali >>
rect -2650 209 -2554 243
rect 2554 209 2650 243
rect -2650 -209 -2616 209
rect -2490 107 -2474 141
rect -2106 107 -2090 141
rect -2032 107 -2016 141
rect -1648 107 -1632 141
rect -1574 107 -1558 141
rect -1190 107 -1174 141
rect -1116 107 -1100 141
rect -732 107 -716 141
rect -658 107 -642 141
rect -274 107 -258 141
rect -200 107 -184 141
rect 184 107 200 141
rect 258 107 274 141
rect 642 107 658 141
rect 716 107 732 141
rect 1100 107 1116 141
rect 1174 107 1190 141
rect 1558 107 1574 141
rect 1632 107 1648 141
rect 2016 107 2032 141
rect 2090 107 2106 141
rect 2474 107 2490 141
rect -2536 57 -2502 73
rect -2536 -135 -2502 -119
rect -2078 57 -2044 73
rect -2078 -135 -2044 -119
rect -1620 57 -1586 73
rect -1620 -135 -1586 -119
rect -1162 57 -1128 73
rect -1162 -135 -1128 -119
rect -704 57 -670 73
rect -704 -135 -670 -119
rect -246 57 -212 73
rect -246 -135 -212 -119
rect 212 57 246 73
rect 212 -135 246 -119
rect 670 57 704 73
rect 670 -135 704 -119
rect 1128 57 1162 73
rect 1128 -135 1162 -119
rect 1586 57 1620 73
rect 1586 -135 1620 -119
rect 2044 57 2078 73
rect 2044 -135 2078 -119
rect 2502 57 2536 73
rect 2502 -135 2536 -119
rect 2616 -209 2650 209
rect -2650 -243 2650 -209
<< viali >>
rect -2474 107 -2106 141
rect -2016 107 -1648 141
rect -1558 107 -1190 141
rect -1100 107 -732 141
rect -642 107 -274 141
rect -184 107 184 141
rect 274 107 642 141
rect 732 107 1100 141
rect 1190 107 1558 141
rect 1648 107 2016 141
rect 2106 107 2474 141
rect -2536 -119 -2502 57
rect -2078 -119 -2044 57
rect -1620 -119 -1586 57
rect -1162 -119 -1128 57
rect -704 -119 -670 57
rect -246 -119 -212 57
rect 212 -119 246 57
rect 670 -119 704 57
rect 1128 -119 1162 57
rect 1586 -119 1620 57
rect 2044 -119 2078 57
rect 2502 -119 2536 57
<< metal1 >>
rect -2486 141 -2094 147
rect -2486 107 -2474 141
rect -2106 107 -2094 141
rect -2486 101 -2094 107
rect -2028 141 -1636 147
rect -2028 107 -2016 141
rect -1648 107 -1636 141
rect -2028 101 -1636 107
rect -1570 141 -1178 147
rect -1570 107 -1558 141
rect -1190 107 -1178 141
rect -1570 101 -1178 107
rect -1112 141 -720 147
rect -1112 107 -1100 141
rect -732 107 -720 141
rect -1112 101 -720 107
rect -654 141 -262 147
rect -654 107 -642 141
rect -274 107 -262 141
rect -654 101 -262 107
rect -196 141 196 147
rect -196 107 -184 141
rect 184 107 196 141
rect -196 101 196 107
rect 262 141 654 147
rect 262 107 274 141
rect 642 107 654 141
rect 262 101 654 107
rect 720 141 1112 147
rect 720 107 732 141
rect 1100 107 1112 141
rect 720 101 1112 107
rect 1178 141 1570 147
rect 1178 107 1190 141
rect 1558 107 1570 141
rect 1178 101 1570 107
rect 1636 141 2028 147
rect 1636 107 1648 141
rect 2016 107 2028 141
rect 1636 101 2028 107
rect 2094 141 2486 147
rect 2094 107 2106 141
rect 2474 107 2486 141
rect 2094 101 2486 107
rect -2542 57 -2496 69
rect -2542 -119 -2536 57
rect -2502 -119 -2496 57
rect -2542 -131 -2496 -119
rect -2084 57 -2038 69
rect -2084 -119 -2078 57
rect -2044 -119 -2038 57
rect -2084 -131 -2038 -119
rect -1626 57 -1580 69
rect -1626 -119 -1620 57
rect -1586 -119 -1580 57
rect -1626 -131 -1580 -119
rect -1168 57 -1122 69
rect -1168 -119 -1162 57
rect -1128 -119 -1122 57
rect -1168 -131 -1122 -119
rect -710 57 -664 69
rect -710 -119 -704 57
rect -670 -119 -664 57
rect -710 -131 -664 -119
rect -252 57 -206 69
rect -252 -119 -246 57
rect -212 -119 -206 57
rect -252 -131 -206 -119
rect 206 57 252 69
rect 206 -119 212 57
rect 246 -119 252 57
rect 206 -131 252 -119
rect 664 57 710 69
rect 664 -119 670 57
rect 704 -119 710 57
rect 664 -131 710 -119
rect 1122 57 1168 69
rect 1122 -119 1128 57
rect 1162 -119 1168 57
rect 1122 -131 1168 -119
rect 1580 57 1626 69
rect 1580 -119 1586 57
rect 1620 -119 1626 57
rect 1580 -131 1626 -119
rect 2038 57 2084 69
rect 2038 -119 2044 57
rect 2078 -119 2084 57
rect 2038 -131 2084 -119
rect 2496 57 2542 69
rect 2496 -119 2502 57
rect 2536 -119 2542 57
rect 2496 -131 2542 -119
<< properties >>
string FIXED_BBOX -2633 -226 2633 226
string gencell sky130_fd_pr__nfet_01v8_lvt
string library sky130
string parameters w 1 l 2 m 1 nf 11 diffcov 100 polycov 100 guard 1 glc 0 grc 0 gtc 1 gbc 0 tbcov 100 rlcov 100 topc 1 botc 0 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
