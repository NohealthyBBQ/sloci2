magic
tech sky130A
magscale 1 2
timestamp 1662761135
<< nwell >>
rect -683 -1014 683 1014
<< pmoslvt >>
rect -487 665 -287 865
rect -229 665 -29 865
rect 29 665 229 865
rect 287 665 487 865
rect -487 300 -287 500
rect -229 300 -29 500
rect 29 300 229 500
rect 287 300 487 500
rect -487 -65 -287 135
rect -229 -65 -29 135
rect 29 -65 229 135
rect 287 -65 487 135
rect -487 -430 -287 -230
rect -229 -430 -29 -230
rect 29 -430 229 -230
rect 287 -430 487 -230
rect -487 -795 -287 -595
rect -229 -795 -29 -595
rect 29 -795 229 -595
rect 287 -795 487 -595
<< pdiff >>
rect -545 853 -487 865
rect -545 677 -533 853
rect -499 677 -487 853
rect -545 665 -487 677
rect -287 853 -229 865
rect -287 677 -275 853
rect -241 677 -229 853
rect -287 665 -229 677
rect -29 853 29 865
rect -29 677 -17 853
rect 17 677 29 853
rect -29 665 29 677
rect 229 853 287 865
rect 229 677 241 853
rect 275 677 287 853
rect 229 665 287 677
rect 487 853 545 865
rect 487 677 499 853
rect 533 677 545 853
rect 487 665 545 677
rect -545 488 -487 500
rect -545 312 -533 488
rect -499 312 -487 488
rect -545 300 -487 312
rect -287 488 -229 500
rect -287 312 -275 488
rect -241 312 -229 488
rect -287 300 -229 312
rect -29 488 29 500
rect -29 312 -17 488
rect 17 312 29 488
rect -29 300 29 312
rect 229 488 287 500
rect 229 312 241 488
rect 275 312 287 488
rect 229 300 287 312
rect 487 488 545 500
rect 487 312 499 488
rect 533 312 545 488
rect 487 300 545 312
rect -545 123 -487 135
rect -545 -53 -533 123
rect -499 -53 -487 123
rect -545 -65 -487 -53
rect -287 123 -229 135
rect -287 -53 -275 123
rect -241 -53 -229 123
rect -287 -65 -229 -53
rect -29 123 29 135
rect -29 -53 -17 123
rect 17 -53 29 123
rect -29 -65 29 -53
rect 229 123 287 135
rect 229 -53 241 123
rect 275 -53 287 123
rect 229 -65 287 -53
rect 487 123 545 135
rect 487 -53 499 123
rect 533 -53 545 123
rect 487 -65 545 -53
rect -545 -242 -487 -230
rect -545 -418 -533 -242
rect -499 -418 -487 -242
rect -545 -430 -487 -418
rect -287 -242 -229 -230
rect -287 -418 -275 -242
rect -241 -418 -229 -242
rect -287 -430 -229 -418
rect -29 -242 29 -230
rect -29 -418 -17 -242
rect 17 -418 29 -242
rect -29 -430 29 -418
rect 229 -242 287 -230
rect 229 -418 241 -242
rect 275 -418 287 -242
rect 229 -430 287 -418
rect 487 -242 545 -230
rect 487 -418 499 -242
rect 533 -418 545 -242
rect 487 -430 545 -418
rect -545 -607 -487 -595
rect -545 -783 -533 -607
rect -499 -783 -487 -607
rect -545 -795 -487 -783
rect -287 -607 -229 -595
rect -287 -783 -275 -607
rect -241 -783 -229 -607
rect -287 -795 -229 -783
rect -29 -607 29 -595
rect -29 -783 -17 -607
rect 17 -783 29 -607
rect -29 -795 29 -783
rect 229 -607 287 -595
rect 229 -783 241 -607
rect 275 -783 287 -607
rect 229 -795 287 -783
rect 487 -607 545 -595
rect 487 -783 499 -607
rect 533 -783 545 -607
rect 487 -795 545 -783
<< pdiffc >>
rect -533 677 -499 853
rect -275 677 -241 853
rect -17 677 17 853
rect 241 677 275 853
rect 499 677 533 853
rect -533 312 -499 488
rect -275 312 -241 488
rect -17 312 17 488
rect 241 312 275 488
rect 499 312 533 488
rect -533 -53 -499 123
rect -275 -53 -241 123
rect -17 -53 17 123
rect 241 -53 275 123
rect 499 -53 533 123
rect -533 -418 -499 -242
rect -275 -418 -241 -242
rect -17 -418 17 -242
rect 241 -418 275 -242
rect 499 -418 533 -242
rect -533 -783 -499 -607
rect -275 -783 -241 -607
rect -17 -783 17 -607
rect 241 -783 275 -607
rect 499 -783 533 -607
<< nsubdiff >>
rect -647 944 -551 978
rect 551 944 647 978
rect -647 882 -613 944
rect 613 882 647 944
rect -647 -944 -613 -882
rect 613 -944 647 -882
rect -647 -978 -551 -944
rect 551 -978 647 -944
<< nsubdiffcont >>
rect -551 944 551 978
rect -647 -882 -613 882
rect 613 -882 647 882
rect -551 -978 551 -944
<< poly >>
rect -487 865 -287 891
rect -229 865 -29 891
rect 29 865 229 891
rect 287 865 487 891
rect -487 618 -287 665
rect -487 584 -471 618
rect -303 584 -287 618
rect -487 568 -287 584
rect -229 618 -29 665
rect -229 584 -213 618
rect -45 584 -29 618
rect -229 568 -29 584
rect 29 618 229 665
rect 29 584 45 618
rect 213 584 229 618
rect 29 568 229 584
rect 287 618 487 665
rect 287 584 303 618
rect 471 584 487 618
rect 287 568 487 584
rect -487 500 -287 526
rect -229 500 -29 526
rect 29 500 229 526
rect 287 500 487 526
rect -487 253 -287 300
rect -487 219 -471 253
rect -303 219 -287 253
rect -487 203 -287 219
rect -229 253 -29 300
rect -229 219 -213 253
rect -45 219 -29 253
rect -229 203 -29 219
rect 29 253 229 300
rect 29 219 45 253
rect 213 219 229 253
rect 29 203 229 219
rect 287 253 487 300
rect 287 219 303 253
rect 471 219 487 253
rect 287 203 487 219
rect -487 135 -287 161
rect -229 135 -29 161
rect 29 135 229 161
rect 287 135 487 161
rect -487 -112 -287 -65
rect -487 -146 -471 -112
rect -303 -146 -287 -112
rect -487 -162 -287 -146
rect -229 -112 -29 -65
rect -229 -146 -213 -112
rect -45 -146 -29 -112
rect -229 -162 -29 -146
rect 29 -112 229 -65
rect 29 -146 45 -112
rect 213 -146 229 -112
rect 29 -162 229 -146
rect 287 -112 487 -65
rect 287 -146 303 -112
rect 471 -146 487 -112
rect 287 -162 487 -146
rect -487 -230 -287 -204
rect -229 -230 -29 -204
rect 29 -230 229 -204
rect 287 -230 487 -204
rect -487 -477 -287 -430
rect -487 -511 -471 -477
rect -303 -511 -287 -477
rect -487 -527 -287 -511
rect -229 -477 -29 -430
rect -229 -511 -213 -477
rect -45 -511 -29 -477
rect -229 -527 -29 -511
rect 29 -477 229 -430
rect 29 -511 45 -477
rect 213 -511 229 -477
rect 29 -527 229 -511
rect 287 -477 487 -430
rect 287 -511 303 -477
rect 471 -511 487 -477
rect 287 -527 487 -511
rect -487 -595 -287 -569
rect -229 -595 -29 -569
rect 29 -595 229 -569
rect 287 -595 487 -569
rect -487 -842 -287 -795
rect -487 -876 -471 -842
rect -303 -876 -287 -842
rect -487 -892 -287 -876
rect -229 -842 -29 -795
rect -229 -876 -213 -842
rect -45 -876 -29 -842
rect -229 -892 -29 -876
rect 29 -842 229 -795
rect 29 -876 45 -842
rect 213 -876 229 -842
rect 29 -892 229 -876
rect 287 -842 487 -795
rect 287 -876 303 -842
rect 471 -876 487 -842
rect 287 -892 487 -876
<< polycont >>
rect -471 584 -303 618
rect -213 584 -45 618
rect 45 584 213 618
rect 303 584 471 618
rect -471 219 -303 253
rect -213 219 -45 253
rect 45 219 213 253
rect 303 219 471 253
rect -471 -146 -303 -112
rect -213 -146 -45 -112
rect 45 -146 213 -112
rect 303 -146 471 -112
rect -471 -511 -303 -477
rect -213 -511 -45 -477
rect 45 -511 213 -477
rect 303 -511 471 -477
rect -471 -876 -303 -842
rect -213 -876 -45 -842
rect 45 -876 213 -842
rect 303 -876 471 -842
<< locali >>
rect -647 944 -551 978
rect 551 944 647 978
rect -647 882 -613 944
rect 613 882 647 944
rect -533 853 -499 869
rect -533 661 -499 677
rect -275 853 -241 869
rect -275 661 -241 677
rect -17 853 17 869
rect -17 661 17 677
rect 241 853 275 869
rect 241 661 275 677
rect 499 853 533 869
rect 499 661 533 677
rect -487 584 -471 618
rect -303 584 -287 618
rect -229 584 -213 618
rect -45 584 -29 618
rect 29 584 45 618
rect 213 584 229 618
rect 287 584 303 618
rect 471 584 487 618
rect -533 488 -499 504
rect -533 296 -499 312
rect -275 488 -241 504
rect -275 296 -241 312
rect -17 488 17 504
rect -17 296 17 312
rect 241 488 275 504
rect 241 296 275 312
rect 499 488 533 504
rect 499 296 533 312
rect -487 219 -471 253
rect -303 219 -287 253
rect -229 219 -213 253
rect -45 219 -29 253
rect 29 219 45 253
rect 213 219 229 253
rect 287 219 303 253
rect 471 219 487 253
rect -533 123 -499 139
rect -533 -69 -499 -53
rect -275 123 -241 139
rect -275 -69 -241 -53
rect -17 123 17 139
rect -17 -69 17 -53
rect 241 123 275 139
rect 241 -69 275 -53
rect 499 123 533 139
rect 499 -69 533 -53
rect -487 -146 -471 -112
rect -303 -146 -287 -112
rect -229 -146 -213 -112
rect -45 -146 -29 -112
rect 29 -146 45 -112
rect 213 -146 229 -112
rect 287 -146 303 -112
rect 471 -146 487 -112
rect -533 -242 -499 -226
rect -533 -434 -499 -418
rect -275 -242 -241 -226
rect -275 -434 -241 -418
rect -17 -242 17 -226
rect -17 -434 17 -418
rect 241 -242 275 -226
rect 241 -434 275 -418
rect 499 -242 533 -226
rect 499 -434 533 -418
rect -487 -511 -471 -477
rect -303 -511 -287 -477
rect -229 -511 -213 -477
rect -45 -511 -29 -477
rect 29 -511 45 -477
rect 213 -511 229 -477
rect 287 -511 303 -477
rect 471 -511 487 -477
rect -533 -607 -499 -591
rect -533 -799 -499 -783
rect -275 -607 -241 -591
rect -275 -799 -241 -783
rect -17 -607 17 -591
rect -17 -799 17 -783
rect 241 -607 275 -591
rect 241 -799 275 -783
rect 499 -607 533 -591
rect 499 -799 533 -783
rect -487 -876 -471 -842
rect -303 -876 -287 -842
rect -229 -876 -213 -842
rect -45 -876 -29 -842
rect 29 -876 45 -842
rect 213 -876 229 -842
rect 287 -876 303 -842
rect 471 -876 487 -842
rect -647 -944 -613 -882
rect 613 -944 647 -882
rect -647 -978 -551 -944
rect 551 -978 647 -944
<< viali >>
rect -533 677 -499 853
rect -275 677 -241 853
rect -17 677 17 853
rect 241 677 275 853
rect 499 677 533 853
rect -471 584 -303 618
rect -213 584 -45 618
rect 45 584 213 618
rect 303 584 471 618
rect -533 312 -499 488
rect -275 312 -241 488
rect -17 312 17 488
rect 241 312 275 488
rect 499 312 533 488
rect -471 219 -303 253
rect -213 219 -45 253
rect 45 219 213 253
rect 303 219 471 253
rect -533 -53 -499 123
rect -275 -53 -241 123
rect -17 -53 17 123
rect 241 -53 275 123
rect 499 -53 533 123
rect -471 -146 -303 -112
rect -213 -146 -45 -112
rect 45 -146 213 -112
rect 303 -146 471 -112
rect -533 -418 -499 -242
rect -275 -418 -241 -242
rect -17 -418 17 -242
rect 241 -418 275 -242
rect 499 -418 533 -242
rect -471 -511 -303 -477
rect -213 -511 -45 -477
rect 45 -511 213 -477
rect 303 -511 471 -477
rect -533 -783 -499 -607
rect -275 -783 -241 -607
rect -17 -783 17 -607
rect 241 -783 275 -607
rect 499 -783 533 -607
rect -471 -876 -303 -842
rect -213 -876 -45 -842
rect 45 -876 213 -842
rect 303 -876 471 -842
<< metal1 >>
rect -539 853 -493 865
rect -539 677 -533 853
rect -499 677 -493 853
rect -539 665 -493 677
rect -281 853 -235 865
rect -281 677 -275 853
rect -241 677 -235 853
rect -281 665 -235 677
rect -23 853 23 865
rect -23 677 -17 853
rect 17 677 23 853
rect -23 665 23 677
rect 235 853 281 865
rect 235 677 241 853
rect 275 677 281 853
rect 235 665 281 677
rect 493 853 539 865
rect 493 677 499 853
rect 533 677 539 853
rect 493 665 539 677
rect -483 618 -291 624
rect -483 584 -471 618
rect -303 584 -291 618
rect -483 578 -291 584
rect -225 618 -33 624
rect -225 584 -213 618
rect -45 584 -33 618
rect -225 578 -33 584
rect 33 618 225 624
rect 33 584 45 618
rect 213 584 225 618
rect 33 578 225 584
rect 291 618 483 624
rect 291 584 303 618
rect 471 584 483 618
rect 291 578 483 584
rect -539 488 -493 500
rect -539 312 -533 488
rect -499 312 -493 488
rect -539 300 -493 312
rect -281 488 -235 500
rect -281 312 -275 488
rect -241 312 -235 488
rect -281 300 -235 312
rect -23 488 23 500
rect -23 312 -17 488
rect 17 312 23 488
rect -23 300 23 312
rect 235 488 281 500
rect 235 312 241 488
rect 275 312 281 488
rect 235 300 281 312
rect 493 488 539 500
rect 493 312 499 488
rect 533 312 539 488
rect 493 300 539 312
rect -483 253 -291 259
rect -483 219 -471 253
rect -303 219 -291 253
rect -483 213 -291 219
rect -225 253 -33 259
rect -225 219 -213 253
rect -45 219 -33 253
rect -225 213 -33 219
rect 33 253 225 259
rect 33 219 45 253
rect 213 219 225 253
rect 33 213 225 219
rect 291 253 483 259
rect 291 219 303 253
rect 471 219 483 253
rect 291 213 483 219
rect -539 123 -493 135
rect -539 -53 -533 123
rect -499 -53 -493 123
rect -539 -65 -493 -53
rect -281 123 -235 135
rect -281 -53 -275 123
rect -241 -53 -235 123
rect -281 -65 -235 -53
rect -23 123 23 135
rect -23 -53 -17 123
rect 17 -53 23 123
rect -23 -65 23 -53
rect 235 123 281 135
rect 235 -53 241 123
rect 275 -53 281 123
rect 235 -65 281 -53
rect 493 123 539 135
rect 493 -53 499 123
rect 533 -53 539 123
rect 493 -65 539 -53
rect -483 -112 -291 -106
rect -483 -146 -471 -112
rect -303 -146 -291 -112
rect -483 -152 -291 -146
rect -225 -112 -33 -106
rect -225 -146 -213 -112
rect -45 -146 -33 -112
rect -225 -152 -33 -146
rect 33 -112 225 -106
rect 33 -146 45 -112
rect 213 -146 225 -112
rect 33 -152 225 -146
rect 291 -112 483 -106
rect 291 -146 303 -112
rect 471 -146 483 -112
rect 291 -152 483 -146
rect -539 -242 -493 -230
rect -539 -418 -533 -242
rect -499 -418 -493 -242
rect -539 -430 -493 -418
rect -281 -242 -235 -230
rect -281 -418 -275 -242
rect -241 -418 -235 -242
rect -281 -430 -235 -418
rect -23 -242 23 -230
rect -23 -418 -17 -242
rect 17 -418 23 -242
rect -23 -430 23 -418
rect 235 -242 281 -230
rect 235 -418 241 -242
rect 275 -418 281 -242
rect 235 -430 281 -418
rect 493 -242 539 -230
rect 493 -418 499 -242
rect 533 -418 539 -242
rect 493 -430 539 -418
rect -483 -477 -291 -471
rect -483 -511 -471 -477
rect -303 -511 -291 -477
rect -483 -517 -291 -511
rect -225 -477 -33 -471
rect -225 -511 -213 -477
rect -45 -511 -33 -477
rect -225 -517 -33 -511
rect 33 -477 225 -471
rect 33 -511 45 -477
rect 213 -511 225 -477
rect 33 -517 225 -511
rect 291 -477 483 -471
rect 291 -511 303 -477
rect 471 -511 483 -477
rect 291 -517 483 -511
rect -539 -607 -493 -595
rect -539 -783 -533 -607
rect -499 -783 -493 -607
rect -539 -795 -493 -783
rect -281 -607 -235 -595
rect -281 -783 -275 -607
rect -241 -783 -235 -607
rect -281 -795 -235 -783
rect -23 -607 23 -595
rect -23 -783 -17 -607
rect 17 -783 23 -607
rect -23 -795 23 -783
rect 235 -607 281 -595
rect 235 -783 241 -607
rect 275 -783 281 -607
rect 235 -795 281 -783
rect 493 -607 539 -595
rect 493 -783 499 -607
rect 533 -783 539 -607
rect 493 -795 539 -783
rect -483 -842 -291 -836
rect -483 -876 -471 -842
rect -303 -876 -291 -842
rect -483 -882 -291 -876
rect -225 -842 -33 -836
rect -225 -876 -213 -842
rect -45 -876 -33 -842
rect -225 -882 -33 -876
rect 33 -842 225 -836
rect 33 -876 45 -842
rect 213 -876 225 -842
rect 33 -882 225 -876
rect 291 -842 483 -836
rect 291 -876 303 -842
rect 471 -876 483 -842
rect 291 -882 483 -876
<< properties >>
string FIXED_BBOX -630 -961 630 961
string gencell sky130_fd_pr__pfet_01v8_lvt
string library sky130
string parameters w 1 l 1 m 5 nf 4 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 0 botc 1 poverlap 0 doverlap 1 lmin 0.35 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
