magic
tech sky130A
magscale 1 2
timestamp 1662478139
<< pwell >>
rect -739 -1190 739 1190
<< psubdiff >>
rect -703 1120 -607 1154
rect 607 1120 703 1154
rect -703 1058 -669 1120
rect 669 1058 703 1120
rect -703 -1120 -669 -1058
rect 669 -1120 703 -1058
rect -703 -1154 -607 -1120
rect 607 -1154 703 -1120
<< psubdiffcont >>
rect -607 1120 607 1154
rect -703 -1058 -669 1058
rect 669 -1058 703 1058
rect -607 -1154 607 -1120
<< xpolycontact >>
rect -573 592 573 1024
rect -573 -1024 573 -592
<< xpolyres >>
rect -573 -592 573 592
<< locali >>
rect -703 1120 -607 1154
rect 607 1120 703 1154
rect -703 1058 -669 1120
rect 669 1058 703 1120
rect -703 -1120 -669 -1058
rect 669 -1120 703 -1058
rect -703 -1154 -607 -1120
rect 607 -1154 703 -1120
<< viali >>
rect -557 609 557 1006
rect -557 -1006 557 -609
<< metal1 >>
rect -569 1006 569 1012
rect -569 609 -557 1006
rect 557 609 569 1006
rect -569 603 569 609
rect -569 -609 569 -603
rect -569 -1006 -557 -609
rect 557 -1006 569 -609
rect -569 -1012 569 -1006
<< res5p73 >>
rect -575 -594 575 594
<< properties >>
string FIXED_BBOX -686 -1137 686 1137
string gencell sky130_fd_pr__res_xhigh_po_5p73
string library sky130
string parameters w 5.730 l 5.92 m 1 nx 1 wmin 5.730 lmin 0.50 rho 2000 val 2.132k dummy 0 dw 0.0 term 188.2 sterm 0.0 caplen 0 wmax 5.730 guard 1 glc 1 grc 1 gtc 1 gbc 1 compatible {sky130_fd_pr__res_xhigh_po_0p35  sky130_fd_pr__res_xhigh_po_0p69 sky130_fd_pr__res_xhigh_po_1p41  sky130_fd_pr__res_xhigh_po_2p85 sky130_fd_pr__res_xhigh_po_5p73} full_metal 1 n_guard 0 hv_guard 0 vias 1 viagb 0 viagt 0 viagl 0 viagr 0
<< end >>
