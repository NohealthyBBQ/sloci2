magic
tech sky130A
magscale 1 2
timestamp 1671758665
<< nwell >>
rect -1747 -1019 1747 1019
<< pmoslvt >>
rect -1551 -800 -1451 800
rect -1393 -800 -1293 800
rect -1235 -800 -1135 800
rect -1077 -800 -977 800
rect -919 -800 -819 800
rect -761 -800 -661 800
rect -603 -800 -503 800
rect -445 -800 -345 800
rect -287 -800 -187 800
rect -129 -800 -29 800
rect 29 -800 129 800
rect 187 -800 287 800
rect 345 -800 445 800
rect 503 -800 603 800
rect 661 -800 761 800
rect 819 -800 919 800
rect 977 -800 1077 800
rect 1135 -800 1235 800
rect 1293 -800 1393 800
rect 1451 -800 1551 800
<< pdiff >>
rect -1609 788 -1551 800
rect -1609 -788 -1597 788
rect -1563 -788 -1551 788
rect -1609 -800 -1551 -788
rect -1451 788 -1393 800
rect -1451 -788 -1439 788
rect -1405 -788 -1393 788
rect -1451 -800 -1393 -788
rect -1293 788 -1235 800
rect -1293 -788 -1281 788
rect -1247 -788 -1235 788
rect -1293 -800 -1235 -788
rect -1135 788 -1077 800
rect -1135 -788 -1123 788
rect -1089 -788 -1077 788
rect -1135 -800 -1077 -788
rect -977 788 -919 800
rect -977 -788 -965 788
rect -931 -788 -919 788
rect -977 -800 -919 -788
rect -819 788 -761 800
rect -819 -788 -807 788
rect -773 -788 -761 788
rect -819 -800 -761 -788
rect -661 788 -603 800
rect -661 -788 -649 788
rect -615 -788 -603 788
rect -661 -800 -603 -788
rect -503 788 -445 800
rect -503 -788 -491 788
rect -457 -788 -445 788
rect -503 -800 -445 -788
rect -345 788 -287 800
rect -345 -788 -333 788
rect -299 -788 -287 788
rect -345 -800 -287 -788
rect -187 788 -129 800
rect -187 -788 -175 788
rect -141 -788 -129 788
rect -187 -800 -129 -788
rect -29 788 29 800
rect -29 -788 -17 788
rect 17 -788 29 788
rect -29 -800 29 -788
rect 129 788 187 800
rect 129 -788 141 788
rect 175 -788 187 788
rect 129 -800 187 -788
rect 287 788 345 800
rect 287 -788 299 788
rect 333 -788 345 788
rect 287 -800 345 -788
rect 445 788 503 800
rect 445 -788 457 788
rect 491 -788 503 788
rect 445 -800 503 -788
rect 603 788 661 800
rect 603 -788 615 788
rect 649 -788 661 788
rect 603 -800 661 -788
rect 761 788 819 800
rect 761 -788 773 788
rect 807 -788 819 788
rect 761 -800 819 -788
rect 919 788 977 800
rect 919 -788 931 788
rect 965 -788 977 788
rect 919 -800 977 -788
rect 1077 788 1135 800
rect 1077 -788 1089 788
rect 1123 -788 1135 788
rect 1077 -800 1135 -788
rect 1235 788 1293 800
rect 1235 -788 1247 788
rect 1281 -788 1293 788
rect 1235 -800 1293 -788
rect 1393 788 1451 800
rect 1393 -788 1405 788
rect 1439 -788 1451 788
rect 1393 -800 1451 -788
rect 1551 788 1609 800
rect 1551 -788 1563 788
rect 1597 -788 1609 788
rect 1551 -800 1609 -788
<< pdiffc >>
rect -1597 -788 -1563 788
rect -1439 -788 -1405 788
rect -1281 -788 -1247 788
rect -1123 -788 -1089 788
rect -965 -788 -931 788
rect -807 -788 -773 788
rect -649 -788 -615 788
rect -491 -788 -457 788
rect -333 -788 -299 788
rect -175 -788 -141 788
rect -17 -788 17 788
rect 141 -788 175 788
rect 299 -788 333 788
rect 457 -788 491 788
rect 615 -788 649 788
rect 773 -788 807 788
rect 931 -788 965 788
rect 1089 -788 1123 788
rect 1247 -788 1281 788
rect 1405 -788 1439 788
rect 1563 -788 1597 788
<< nsubdiff >>
rect -1711 949 -1615 983
rect 1615 949 1711 983
rect -1711 -949 -1677 949
rect 1677 -949 1711 949
rect -1711 -983 -1615 -949
rect 1615 -983 1711 -949
<< nsubdiffcont >>
rect -1615 949 1615 983
rect -1615 -983 1615 -949
<< poly >>
rect -1551 881 -1451 897
rect -1551 847 -1535 881
rect -1467 847 -1451 881
rect -1551 800 -1451 847
rect -1393 881 -1293 897
rect -1393 847 -1377 881
rect -1309 847 -1293 881
rect -1393 800 -1293 847
rect -1235 881 -1135 897
rect -1235 847 -1219 881
rect -1151 847 -1135 881
rect -1235 800 -1135 847
rect -1077 881 -977 897
rect -1077 847 -1061 881
rect -993 847 -977 881
rect -1077 800 -977 847
rect -919 881 -819 897
rect -919 847 -903 881
rect -835 847 -819 881
rect -919 800 -819 847
rect -761 881 -661 897
rect -761 847 -745 881
rect -677 847 -661 881
rect -761 800 -661 847
rect -603 881 -503 897
rect -603 847 -587 881
rect -519 847 -503 881
rect -603 800 -503 847
rect -445 881 -345 897
rect -445 847 -429 881
rect -361 847 -345 881
rect -445 800 -345 847
rect -287 881 -187 897
rect -287 847 -271 881
rect -203 847 -187 881
rect -287 800 -187 847
rect -129 881 -29 897
rect -129 847 -113 881
rect -45 847 -29 881
rect -129 800 -29 847
rect 29 881 129 897
rect 29 847 45 881
rect 113 847 129 881
rect 29 800 129 847
rect 187 881 287 897
rect 187 847 203 881
rect 271 847 287 881
rect 187 800 287 847
rect 345 881 445 897
rect 345 847 361 881
rect 429 847 445 881
rect 345 800 445 847
rect 503 881 603 897
rect 503 847 519 881
rect 587 847 603 881
rect 503 800 603 847
rect 661 881 761 897
rect 661 847 677 881
rect 745 847 761 881
rect 661 800 761 847
rect 819 881 919 897
rect 819 847 835 881
rect 903 847 919 881
rect 819 800 919 847
rect 977 881 1077 897
rect 977 847 993 881
rect 1061 847 1077 881
rect 977 800 1077 847
rect 1135 881 1235 897
rect 1135 847 1151 881
rect 1219 847 1235 881
rect 1135 800 1235 847
rect 1293 881 1393 897
rect 1293 847 1309 881
rect 1377 847 1393 881
rect 1293 800 1393 847
rect 1451 881 1551 897
rect 1451 847 1467 881
rect 1535 847 1551 881
rect 1451 800 1551 847
rect -1551 -847 -1451 -800
rect -1551 -881 -1535 -847
rect -1467 -881 -1451 -847
rect -1551 -897 -1451 -881
rect -1393 -847 -1293 -800
rect -1393 -881 -1377 -847
rect -1309 -881 -1293 -847
rect -1393 -897 -1293 -881
rect -1235 -847 -1135 -800
rect -1235 -881 -1219 -847
rect -1151 -881 -1135 -847
rect -1235 -897 -1135 -881
rect -1077 -847 -977 -800
rect -1077 -881 -1061 -847
rect -993 -881 -977 -847
rect -1077 -897 -977 -881
rect -919 -847 -819 -800
rect -919 -881 -903 -847
rect -835 -881 -819 -847
rect -919 -897 -819 -881
rect -761 -847 -661 -800
rect -761 -881 -745 -847
rect -677 -881 -661 -847
rect -761 -897 -661 -881
rect -603 -847 -503 -800
rect -603 -881 -587 -847
rect -519 -881 -503 -847
rect -603 -897 -503 -881
rect -445 -847 -345 -800
rect -445 -881 -429 -847
rect -361 -881 -345 -847
rect -445 -897 -345 -881
rect -287 -847 -187 -800
rect -287 -881 -271 -847
rect -203 -881 -187 -847
rect -287 -897 -187 -881
rect -129 -847 -29 -800
rect -129 -881 -113 -847
rect -45 -881 -29 -847
rect -129 -897 -29 -881
rect 29 -847 129 -800
rect 29 -881 45 -847
rect 113 -881 129 -847
rect 29 -897 129 -881
rect 187 -847 287 -800
rect 187 -881 203 -847
rect 271 -881 287 -847
rect 187 -897 287 -881
rect 345 -847 445 -800
rect 345 -881 361 -847
rect 429 -881 445 -847
rect 345 -897 445 -881
rect 503 -847 603 -800
rect 503 -881 519 -847
rect 587 -881 603 -847
rect 503 -897 603 -881
rect 661 -847 761 -800
rect 661 -881 677 -847
rect 745 -881 761 -847
rect 661 -897 761 -881
rect 819 -847 919 -800
rect 819 -881 835 -847
rect 903 -881 919 -847
rect 819 -897 919 -881
rect 977 -847 1077 -800
rect 977 -881 993 -847
rect 1061 -881 1077 -847
rect 977 -897 1077 -881
rect 1135 -847 1235 -800
rect 1135 -881 1151 -847
rect 1219 -881 1235 -847
rect 1135 -897 1235 -881
rect 1293 -847 1393 -800
rect 1293 -881 1309 -847
rect 1377 -881 1393 -847
rect 1293 -897 1393 -881
rect 1451 -847 1551 -800
rect 1451 -881 1467 -847
rect 1535 -881 1551 -847
rect 1451 -897 1551 -881
<< polycont >>
rect -1535 847 -1467 881
rect -1377 847 -1309 881
rect -1219 847 -1151 881
rect -1061 847 -993 881
rect -903 847 -835 881
rect -745 847 -677 881
rect -587 847 -519 881
rect -429 847 -361 881
rect -271 847 -203 881
rect -113 847 -45 881
rect 45 847 113 881
rect 203 847 271 881
rect 361 847 429 881
rect 519 847 587 881
rect 677 847 745 881
rect 835 847 903 881
rect 993 847 1061 881
rect 1151 847 1219 881
rect 1309 847 1377 881
rect 1467 847 1535 881
rect -1535 -881 -1467 -847
rect -1377 -881 -1309 -847
rect -1219 -881 -1151 -847
rect -1061 -881 -993 -847
rect -903 -881 -835 -847
rect -745 -881 -677 -847
rect -587 -881 -519 -847
rect -429 -881 -361 -847
rect -271 -881 -203 -847
rect -113 -881 -45 -847
rect 45 -881 113 -847
rect 203 -881 271 -847
rect 361 -881 429 -847
rect 519 -881 587 -847
rect 677 -881 745 -847
rect 835 -881 903 -847
rect 993 -881 1061 -847
rect 1151 -881 1219 -847
rect 1309 -881 1377 -847
rect 1467 -881 1535 -847
<< locali >>
rect -1711 949 -1615 983
rect 1615 949 1711 983
rect -1711 -949 -1677 949
rect -1551 847 -1535 881
rect -1467 847 -1451 881
rect -1393 847 -1377 881
rect -1309 847 -1293 881
rect -1235 847 -1219 881
rect -1151 847 -1135 881
rect -1077 847 -1061 881
rect -993 847 -977 881
rect -919 847 -903 881
rect -835 847 -819 881
rect -761 847 -745 881
rect -677 847 -661 881
rect -603 847 -587 881
rect -519 847 -503 881
rect -445 847 -429 881
rect -361 847 -345 881
rect -287 847 -271 881
rect -203 847 -187 881
rect -129 847 -113 881
rect -45 847 -29 881
rect 29 847 45 881
rect 113 847 129 881
rect 187 847 203 881
rect 271 847 287 881
rect 345 847 361 881
rect 429 847 445 881
rect 503 847 519 881
rect 587 847 603 881
rect 661 847 677 881
rect 745 847 761 881
rect 819 847 835 881
rect 903 847 919 881
rect 977 847 993 881
rect 1061 847 1077 881
rect 1135 847 1151 881
rect 1219 847 1235 881
rect 1293 847 1309 881
rect 1377 847 1393 881
rect 1451 847 1467 881
rect 1535 847 1551 881
rect -1597 788 -1563 804
rect -1597 -804 -1563 -788
rect -1439 788 -1405 804
rect -1439 -804 -1405 -788
rect -1281 788 -1247 804
rect -1281 -804 -1247 -788
rect -1123 788 -1089 804
rect -1123 -804 -1089 -788
rect -965 788 -931 804
rect -965 -804 -931 -788
rect -807 788 -773 804
rect -807 -804 -773 -788
rect -649 788 -615 804
rect -649 -804 -615 -788
rect -491 788 -457 804
rect -491 -804 -457 -788
rect -333 788 -299 804
rect -333 -804 -299 -788
rect -175 788 -141 804
rect -175 -804 -141 -788
rect -17 788 17 804
rect -17 -804 17 -788
rect 141 788 175 804
rect 141 -804 175 -788
rect 299 788 333 804
rect 299 -804 333 -788
rect 457 788 491 804
rect 457 -804 491 -788
rect 615 788 649 804
rect 615 -804 649 -788
rect 773 788 807 804
rect 773 -804 807 -788
rect 931 788 965 804
rect 931 -804 965 -788
rect 1089 788 1123 804
rect 1089 -804 1123 -788
rect 1247 788 1281 804
rect 1247 -804 1281 -788
rect 1405 788 1439 804
rect 1405 -804 1439 -788
rect 1563 788 1597 804
rect 1563 -804 1597 -788
rect -1551 -881 -1535 -847
rect -1467 -881 -1451 -847
rect -1393 -881 -1377 -847
rect -1309 -881 -1293 -847
rect -1235 -881 -1219 -847
rect -1151 -881 -1135 -847
rect -1077 -881 -1061 -847
rect -993 -881 -977 -847
rect -919 -881 -903 -847
rect -835 -881 -819 -847
rect -761 -881 -745 -847
rect -677 -881 -661 -847
rect -603 -881 -587 -847
rect -519 -881 -503 -847
rect -445 -881 -429 -847
rect -361 -881 -345 -847
rect -287 -881 -271 -847
rect -203 -881 -187 -847
rect -129 -881 -113 -847
rect -45 -881 -29 -847
rect 29 -881 45 -847
rect 113 -881 129 -847
rect 187 -881 203 -847
rect 271 -881 287 -847
rect 345 -881 361 -847
rect 429 -881 445 -847
rect 503 -881 519 -847
rect 587 -881 603 -847
rect 661 -881 677 -847
rect 745 -881 761 -847
rect 819 -881 835 -847
rect 903 -881 919 -847
rect 977 -881 993 -847
rect 1061 -881 1077 -847
rect 1135 -881 1151 -847
rect 1219 -881 1235 -847
rect 1293 -881 1309 -847
rect 1377 -881 1393 -847
rect 1451 -881 1467 -847
rect 1535 -881 1551 -847
rect 1677 -949 1711 949
rect -1711 -983 -1615 -949
rect 1615 -983 1711 -949
<< viali >>
rect -1535 847 -1467 881
rect -1377 847 -1309 881
rect -1219 847 -1151 881
rect -1061 847 -993 881
rect -903 847 -835 881
rect -745 847 -677 881
rect -587 847 -519 881
rect -429 847 -361 881
rect -271 847 -203 881
rect -113 847 -45 881
rect 45 847 113 881
rect 203 847 271 881
rect 361 847 429 881
rect 519 847 587 881
rect 677 847 745 881
rect 835 847 903 881
rect 993 847 1061 881
rect 1151 847 1219 881
rect 1309 847 1377 881
rect 1467 847 1535 881
rect -1597 -788 -1563 788
rect -1439 -788 -1405 788
rect -1281 -788 -1247 788
rect -1123 -788 -1089 788
rect -965 -788 -931 788
rect -807 -788 -773 788
rect -649 -788 -615 788
rect -491 -788 -457 788
rect -333 -788 -299 788
rect -175 -788 -141 788
rect -17 -788 17 788
rect 141 -788 175 788
rect 299 -788 333 788
rect 457 -788 491 788
rect 615 -788 649 788
rect 773 -788 807 788
rect 931 -788 965 788
rect 1089 -788 1123 788
rect 1247 -788 1281 788
rect 1405 -788 1439 788
rect 1563 -788 1597 788
rect -1535 -881 -1467 -847
rect -1377 -881 -1309 -847
rect -1219 -881 -1151 -847
rect -1061 -881 -993 -847
rect -903 -881 -835 -847
rect -745 -881 -677 -847
rect -587 -881 -519 -847
rect -429 -881 -361 -847
rect -271 -881 -203 -847
rect -113 -881 -45 -847
rect 45 -881 113 -847
rect 203 -881 271 -847
rect 361 -881 429 -847
rect 519 -881 587 -847
rect 677 -881 745 -847
rect 835 -881 903 -847
rect 993 -881 1061 -847
rect 1151 -881 1219 -847
rect 1309 -881 1377 -847
rect 1467 -881 1535 -847
<< metal1 >>
rect -1547 881 -1455 887
rect -1547 847 -1535 881
rect -1467 847 -1455 881
rect -1547 841 -1455 847
rect -1389 881 -1297 887
rect -1389 847 -1377 881
rect -1309 847 -1297 881
rect -1389 841 -1297 847
rect -1231 881 -1139 887
rect -1231 847 -1219 881
rect -1151 847 -1139 881
rect -1231 841 -1139 847
rect -1073 881 -981 887
rect -1073 847 -1061 881
rect -993 847 -981 881
rect -1073 841 -981 847
rect -915 881 -823 887
rect -915 847 -903 881
rect -835 847 -823 881
rect -915 841 -823 847
rect -757 881 -665 887
rect -757 847 -745 881
rect -677 847 -665 881
rect -757 841 -665 847
rect -599 881 -507 887
rect -599 847 -587 881
rect -519 847 -507 881
rect -599 841 -507 847
rect -441 881 -349 887
rect -441 847 -429 881
rect -361 847 -349 881
rect -441 841 -349 847
rect -283 881 -191 887
rect -283 847 -271 881
rect -203 847 -191 881
rect -283 841 -191 847
rect -125 881 -33 887
rect -125 847 -113 881
rect -45 847 -33 881
rect -125 841 -33 847
rect 33 881 125 887
rect 33 847 45 881
rect 113 847 125 881
rect 33 841 125 847
rect 191 881 283 887
rect 191 847 203 881
rect 271 847 283 881
rect 191 841 283 847
rect 349 881 441 887
rect 349 847 361 881
rect 429 847 441 881
rect 349 841 441 847
rect 507 881 599 887
rect 507 847 519 881
rect 587 847 599 881
rect 507 841 599 847
rect 665 881 757 887
rect 665 847 677 881
rect 745 847 757 881
rect 665 841 757 847
rect 823 881 915 887
rect 823 847 835 881
rect 903 847 915 881
rect 823 841 915 847
rect 981 881 1073 887
rect 981 847 993 881
rect 1061 847 1073 881
rect 981 841 1073 847
rect 1139 881 1231 887
rect 1139 847 1151 881
rect 1219 847 1231 881
rect 1139 841 1231 847
rect 1297 881 1389 887
rect 1297 847 1309 881
rect 1377 847 1389 881
rect 1297 841 1389 847
rect 1455 881 1547 887
rect 1455 847 1467 881
rect 1535 847 1547 881
rect 1455 841 1547 847
rect -1603 788 -1557 800
rect -1603 -788 -1597 788
rect -1563 -788 -1557 788
rect -1603 -800 -1557 -788
rect -1445 788 -1399 800
rect -1445 -788 -1439 788
rect -1405 -788 -1399 788
rect -1445 -800 -1399 -788
rect -1287 788 -1241 800
rect -1287 -788 -1281 788
rect -1247 -788 -1241 788
rect -1287 -800 -1241 -788
rect -1129 788 -1083 800
rect -1129 -788 -1123 788
rect -1089 -788 -1083 788
rect -1129 -800 -1083 -788
rect -971 788 -925 800
rect -971 -788 -965 788
rect -931 -788 -925 788
rect -971 -800 -925 -788
rect -813 788 -767 800
rect -813 -788 -807 788
rect -773 -788 -767 788
rect -813 -800 -767 -788
rect -655 788 -609 800
rect -655 -788 -649 788
rect -615 -788 -609 788
rect -655 -800 -609 -788
rect -497 788 -451 800
rect -497 -788 -491 788
rect -457 -788 -451 788
rect -497 -800 -451 -788
rect -339 788 -293 800
rect -339 -788 -333 788
rect -299 -788 -293 788
rect -339 -800 -293 -788
rect -181 788 -135 800
rect -181 -788 -175 788
rect -141 -788 -135 788
rect -181 -800 -135 -788
rect -23 788 23 800
rect -23 -788 -17 788
rect 17 -788 23 788
rect -23 -800 23 -788
rect 135 788 181 800
rect 135 -788 141 788
rect 175 -788 181 788
rect 135 -800 181 -788
rect 293 788 339 800
rect 293 -788 299 788
rect 333 -788 339 788
rect 293 -800 339 -788
rect 451 788 497 800
rect 451 -788 457 788
rect 491 -788 497 788
rect 451 -800 497 -788
rect 609 788 655 800
rect 609 -788 615 788
rect 649 -788 655 788
rect 609 -800 655 -788
rect 767 788 813 800
rect 767 -788 773 788
rect 807 -788 813 788
rect 767 -800 813 -788
rect 925 788 971 800
rect 925 -788 931 788
rect 965 -788 971 788
rect 925 -800 971 -788
rect 1083 788 1129 800
rect 1083 -788 1089 788
rect 1123 -788 1129 788
rect 1083 -800 1129 -788
rect 1241 788 1287 800
rect 1241 -788 1247 788
rect 1281 -788 1287 788
rect 1241 -800 1287 -788
rect 1399 788 1445 800
rect 1399 -788 1405 788
rect 1439 -788 1445 788
rect 1399 -800 1445 -788
rect 1557 788 1603 800
rect 1557 -788 1563 788
rect 1597 -788 1603 788
rect 1557 -800 1603 -788
rect -1547 -847 -1455 -841
rect -1547 -881 -1535 -847
rect -1467 -881 -1455 -847
rect -1547 -887 -1455 -881
rect -1389 -847 -1297 -841
rect -1389 -881 -1377 -847
rect -1309 -881 -1297 -847
rect -1389 -887 -1297 -881
rect -1231 -847 -1139 -841
rect -1231 -881 -1219 -847
rect -1151 -881 -1139 -847
rect -1231 -887 -1139 -881
rect -1073 -847 -981 -841
rect -1073 -881 -1061 -847
rect -993 -881 -981 -847
rect -1073 -887 -981 -881
rect -915 -847 -823 -841
rect -915 -881 -903 -847
rect -835 -881 -823 -847
rect -915 -887 -823 -881
rect -757 -847 -665 -841
rect -757 -881 -745 -847
rect -677 -881 -665 -847
rect -757 -887 -665 -881
rect -599 -847 -507 -841
rect -599 -881 -587 -847
rect -519 -881 -507 -847
rect -599 -887 -507 -881
rect -441 -847 -349 -841
rect -441 -881 -429 -847
rect -361 -881 -349 -847
rect -441 -887 -349 -881
rect -283 -847 -191 -841
rect -283 -881 -271 -847
rect -203 -881 -191 -847
rect -283 -887 -191 -881
rect -125 -847 -33 -841
rect -125 -881 -113 -847
rect -45 -881 -33 -847
rect -125 -887 -33 -881
rect 33 -847 125 -841
rect 33 -881 45 -847
rect 113 -881 125 -847
rect 33 -887 125 -881
rect 191 -847 283 -841
rect 191 -881 203 -847
rect 271 -881 283 -847
rect 191 -887 283 -881
rect 349 -847 441 -841
rect 349 -881 361 -847
rect 429 -881 441 -847
rect 349 -887 441 -881
rect 507 -847 599 -841
rect 507 -881 519 -847
rect 587 -881 599 -847
rect 507 -887 599 -881
rect 665 -847 757 -841
rect 665 -881 677 -847
rect 745 -881 757 -847
rect 665 -887 757 -881
rect 823 -847 915 -841
rect 823 -881 835 -847
rect 903 -881 915 -847
rect 823 -887 915 -881
rect 981 -847 1073 -841
rect 981 -881 993 -847
rect 1061 -881 1073 -847
rect 981 -887 1073 -881
rect 1139 -847 1231 -841
rect 1139 -881 1151 -847
rect 1219 -881 1231 -847
rect 1139 -887 1231 -881
rect 1297 -847 1389 -841
rect 1297 -881 1309 -847
rect 1377 -881 1389 -847
rect 1297 -887 1389 -881
rect 1455 -847 1547 -841
rect 1455 -881 1467 -847
rect 1535 -881 1547 -847
rect 1455 -887 1547 -881
<< properties >>
string FIXED_BBOX -1694 -966 1694 966
string gencell sky130_fd_pr__pfet_01v8_lvt
string library sky130
string parameters w 8 l 0.5 m 1 nf 20 diffcov 100 polycov 100 guard 1 glc 0 grc 0 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.35 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
