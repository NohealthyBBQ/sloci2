magic
tech sky130A
magscale 1 2
timestamp 1671758665
<< nwell >>
rect -957 -1937 957 1937
<< pmoslvt >>
rect -761 118 -661 1718
rect -603 118 -503 1718
rect -445 118 -345 1718
rect -287 118 -187 1718
rect -129 118 -29 1718
rect 29 118 129 1718
rect 187 118 287 1718
rect 345 118 445 1718
rect 503 118 603 1718
rect 661 118 761 1718
rect -761 -1718 -661 -118
rect -603 -1718 -503 -118
rect -445 -1718 -345 -118
rect -287 -1718 -187 -118
rect -129 -1718 -29 -118
rect 29 -1718 129 -118
rect 187 -1718 287 -118
rect 345 -1718 445 -118
rect 503 -1718 603 -118
rect 661 -1718 761 -118
<< pdiff >>
rect -819 1706 -761 1718
rect -819 130 -807 1706
rect -773 130 -761 1706
rect -819 118 -761 130
rect -661 1706 -603 1718
rect -661 130 -649 1706
rect -615 130 -603 1706
rect -661 118 -603 130
rect -503 1706 -445 1718
rect -503 130 -491 1706
rect -457 130 -445 1706
rect -503 118 -445 130
rect -345 1706 -287 1718
rect -345 130 -333 1706
rect -299 130 -287 1706
rect -345 118 -287 130
rect -187 1706 -129 1718
rect -187 130 -175 1706
rect -141 130 -129 1706
rect -187 118 -129 130
rect -29 1706 29 1718
rect -29 130 -17 1706
rect 17 130 29 1706
rect -29 118 29 130
rect 129 1706 187 1718
rect 129 130 141 1706
rect 175 130 187 1706
rect 129 118 187 130
rect 287 1706 345 1718
rect 287 130 299 1706
rect 333 130 345 1706
rect 287 118 345 130
rect 445 1706 503 1718
rect 445 130 457 1706
rect 491 130 503 1706
rect 445 118 503 130
rect 603 1706 661 1718
rect 603 130 615 1706
rect 649 130 661 1706
rect 603 118 661 130
rect 761 1706 819 1718
rect 761 130 773 1706
rect 807 130 819 1706
rect 761 118 819 130
rect -819 -130 -761 -118
rect -819 -1706 -807 -130
rect -773 -1706 -761 -130
rect -819 -1718 -761 -1706
rect -661 -130 -603 -118
rect -661 -1706 -649 -130
rect -615 -1706 -603 -130
rect -661 -1718 -603 -1706
rect -503 -130 -445 -118
rect -503 -1706 -491 -130
rect -457 -1706 -445 -130
rect -503 -1718 -445 -1706
rect -345 -130 -287 -118
rect -345 -1706 -333 -130
rect -299 -1706 -287 -130
rect -345 -1718 -287 -1706
rect -187 -130 -129 -118
rect -187 -1706 -175 -130
rect -141 -1706 -129 -130
rect -187 -1718 -129 -1706
rect -29 -130 29 -118
rect -29 -1706 -17 -130
rect 17 -1706 29 -130
rect -29 -1718 29 -1706
rect 129 -130 187 -118
rect 129 -1706 141 -130
rect 175 -1706 187 -130
rect 129 -1718 187 -1706
rect 287 -130 345 -118
rect 287 -1706 299 -130
rect 333 -1706 345 -130
rect 287 -1718 345 -1706
rect 445 -130 503 -118
rect 445 -1706 457 -130
rect 491 -1706 503 -130
rect 445 -1718 503 -1706
rect 603 -130 661 -118
rect 603 -1706 615 -130
rect 649 -1706 661 -130
rect 603 -1718 661 -1706
rect 761 -130 819 -118
rect 761 -1706 773 -130
rect 807 -1706 819 -130
rect 761 -1718 819 -1706
<< pdiffc >>
rect -807 130 -773 1706
rect -649 130 -615 1706
rect -491 130 -457 1706
rect -333 130 -299 1706
rect -175 130 -141 1706
rect -17 130 17 1706
rect 141 130 175 1706
rect 299 130 333 1706
rect 457 130 491 1706
rect 615 130 649 1706
rect 773 130 807 1706
rect -807 -1706 -773 -130
rect -649 -1706 -615 -130
rect -491 -1706 -457 -130
rect -333 -1706 -299 -130
rect -175 -1706 -141 -130
rect -17 -1706 17 -130
rect 141 -1706 175 -130
rect 299 -1706 333 -130
rect 457 -1706 491 -130
rect 615 -1706 649 -130
rect 773 -1706 807 -130
<< nsubdiff >>
rect -921 1867 -825 1901
rect 825 1867 921 1901
rect -921 -1867 -887 1867
rect 887 -1867 921 1867
rect -921 -1901 -825 -1867
rect 825 -1901 921 -1867
<< nsubdiffcont >>
rect -825 1867 825 1901
rect -825 -1901 825 -1867
<< poly >>
rect -761 1799 -661 1815
rect -761 1765 -745 1799
rect -677 1765 -661 1799
rect -761 1718 -661 1765
rect -603 1799 -503 1815
rect -603 1765 -587 1799
rect -519 1765 -503 1799
rect -603 1718 -503 1765
rect -445 1799 -345 1815
rect -445 1765 -429 1799
rect -361 1765 -345 1799
rect -445 1718 -345 1765
rect -287 1799 -187 1815
rect -287 1765 -271 1799
rect -203 1765 -187 1799
rect -287 1718 -187 1765
rect -129 1799 -29 1815
rect -129 1765 -113 1799
rect -45 1765 -29 1799
rect -129 1718 -29 1765
rect 29 1799 129 1815
rect 29 1765 45 1799
rect 113 1765 129 1799
rect 29 1718 129 1765
rect 187 1799 287 1815
rect 187 1765 203 1799
rect 271 1765 287 1799
rect 187 1718 287 1765
rect 345 1799 445 1815
rect 345 1765 361 1799
rect 429 1765 445 1799
rect 345 1718 445 1765
rect 503 1799 603 1815
rect 503 1765 519 1799
rect 587 1765 603 1799
rect 503 1718 603 1765
rect 661 1799 761 1815
rect 661 1765 677 1799
rect 745 1765 761 1799
rect 661 1718 761 1765
rect -761 71 -661 118
rect -761 37 -745 71
rect -677 37 -661 71
rect -761 21 -661 37
rect -603 71 -503 118
rect -603 37 -587 71
rect -519 37 -503 71
rect -603 21 -503 37
rect -445 71 -345 118
rect -445 37 -429 71
rect -361 37 -345 71
rect -445 21 -345 37
rect -287 71 -187 118
rect -287 37 -271 71
rect -203 37 -187 71
rect -287 21 -187 37
rect -129 71 -29 118
rect -129 37 -113 71
rect -45 37 -29 71
rect -129 21 -29 37
rect 29 71 129 118
rect 29 37 45 71
rect 113 37 129 71
rect 29 21 129 37
rect 187 71 287 118
rect 187 37 203 71
rect 271 37 287 71
rect 187 21 287 37
rect 345 71 445 118
rect 345 37 361 71
rect 429 37 445 71
rect 345 21 445 37
rect 503 71 603 118
rect 503 37 519 71
rect 587 37 603 71
rect 503 21 603 37
rect 661 71 761 118
rect 661 37 677 71
rect 745 37 761 71
rect 661 21 761 37
rect -761 -37 -661 -21
rect -761 -71 -745 -37
rect -677 -71 -661 -37
rect -761 -118 -661 -71
rect -603 -37 -503 -21
rect -603 -71 -587 -37
rect -519 -71 -503 -37
rect -603 -118 -503 -71
rect -445 -37 -345 -21
rect -445 -71 -429 -37
rect -361 -71 -345 -37
rect -445 -118 -345 -71
rect -287 -37 -187 -21
rect -287 -71 -271 -37
rect -203 -71 -187 -37
rect -287 -118 -187 -71
rect -129 -37 -29 -21
rect -129 -71 -113 -37
rect -45 -71 -29 -37
rect -129 -118 -29 -71
rect 29 -37 129 -21
rect 29 -71 45 -37
rect 113 -71 129 -37
rect 29 -118 129 -71
rect 187 -37 287 -21
rect 187 -71 203 -37
rect 271 -71 287 -37
rect 187 -118 287 -71
rect 345 -37 445 -21
rect 345 -71 361 -37
rect 429 -71 445 -37
rect 345 -118 445 -71
rect 503 -37 603 -21
rect 503 -71 519 -37
rect 587 -71 603 -37
rect 503 -118 603 -71
rect 661 -37 761 -21
rect 661 -71 677 -37
rect 745 -71 761 -37
rect 661 -118 761 -71
rect -761 -1765 -661 -1718
rect -761 -1799 -745 -1765
rect -677 -1799 -661 -1765
rect -761 -1815 -661 -1799
rect -603 -1765 -503 -1718
rect -603 -1799 -587 -1765
rect -519 -1799 -503 -1765
rect -603 -1815 -503 -1799
rect -445 -1765 -345 -1718
rect -445 -1799 -429 -1765
rect -361 -1799 -345 -1765
rect -445 -1815 -345 -1799
rect -287 -1765 -187 -1718
rect -287 -1799 -271 -1765
rect -203 -1799 -187 -1765
rect -287 -1815 -187 -1799
rect -129 -1765 -29 -1718
rect -129 -1799 -113 -1765
rect -45 -1799 -29 -1765
rect -129 -1815 -29 -1799
rect 29 -1765 129 -1718
rect 29 -1799 45 -1765
rect 113 -1799 129 -1765
rect 29 -1815 129 -1799
rect 187 -1765 287 -1718
rect 187 -1799 203 -1765
rect 271 -1799 287 -1765
rect 187 -1815 287 -1799
rect 345 -1765 445 -1718
rect 345 -1799 361 -1765
rect 429 -1799 445 -1765
rect 345 -1815 445 -1799
rect 503 -1765 603 -1718
rect 503 -1799 519 -1765
rect 587 -1799 603 -1765
rect 503 -1815 603 -1799
rect 661 -1765 761 -1718
rect 661 -1799 677 -1765
rect 745 -1799 761 -1765
rect 661 -1815 761 -1799
<< polycont >>
rect -745 1765 -677 1799
rect -587 1765 -519 1799
rect -429 1765 -361 1799
rect -271 1765 -203 1799
rect -113 1765 -45 1799
rect 45 1765 113 1799
rect 203 1765 271 1799
rect 361 1765 429 1799
rect 519 1765 587 1799
rect 677 1765 745 1799
rect -745 37 -677 71
rect -587 37 -519 71
rect -429 37 -361 71
rect -271 37 -203 71
rect -113 37 -45 71
rect 45 37 113 71
rect 203 37 271 71
rect 361 37 429 71
rect 519 37 587 71
rect 677 37 745 71
rect -745 -71 -677 -37
rect -587 -71 -519 -37
rect -429 -71 -361 -37
rect -271 -71 -203 -37
rect -113 -71 -45 -37
rect 45 -71 113 -37
rect 203 -71 271 -37
rect 361 -71 429 -37
rect 519 -71 587 -37
rect 677 -71 745 -37
rect -745 -1799 -677 -1765
rect -587 -1799 -519 -1765
rect -429 -1799 -361 -1765
rect -271 -1799 -203 -1765
rect -113 -1799 -45 -1765
rect 45 -1799 113 -1765
rect 203 -1799 271 -1765
rect 361 -1799 429 -1765
rect 519 -1799 587 -1765
rect 677 -1799 745 -1765
<< locali >>
rect -921 1867 -825 1901
rect 825 1867 921 1901
rect -921 -1867 -887 1867
rect -761 1765 -745 1799
rect -677 1765 -661 1799
rect -603 1765 -587 1799
rect -519 1765 -503 1799
rect -445 1765 -429 1799
rect -361 1765 -345 1799
rect -287 1765 -271 1799
rect -203 1765 -187 1799
rect -129 1765 -113 1799
rect -45 1765 -29 1799
rect 29 1765 45 1799
rect 113 1765 129 1799
rect 187 1765 203 1799
rect 271 1765 287 1799
rect 345 1765 361 1799
rect 429 1765 445 1799
rect 503 1765 519 1799
rect 587 1765 603 1799
rect 661 1765 677 1799
rect 745 1765 761 1799
rect -807 1706 -773 1722
rect -807 114 -773 130
rect -649 1706 -615 1722
rect -649 114 -615 130
rect -491 1706 -457 1722
rect -491 114 -457 130
rect -333 1706 -299 1722
rect -333 114 -299 130
rect -175 1706 -141 1722
rect -175 114 -141 130
rect -17 1706 17 1722
rect -17 114 17 130
rect 141 1706 175 1722
rect 141 114 175 130
rect 299 1706 333 1722
rect 299 114 333 130
rect 457 1706 491 1722
rect 457 114 491 130
rect 615 1706 649 1722
rect 615 114 649 130
rect 773 1706 807 1722
rect 773 114 807 130
rect -761 37 -745 71
rect -677 37 -661 71
rect -603 37 -587 71
rect -519 37 -503 71
rect -445 37 -429 71
rect -361 37 -345 71
rect -287 37 -271 71
rect -203 37 -187 71
rect -129 37 -113 71
rect -45 37 -29 71
rect 29 37 45 71
rect 113 37 129 71
rect 187 37 203 71
rect 271 37 287 71
rect 345 37 361 71
rect 429 37 445 71
rect 503 37 519 71
rect 587 37 603 71
rect 661 37 677 71
rect 745 37 761 71
rect -761 -71 -745 -37
rect -677 -71 -661 -37
rect -603 -71 -587 -37
rect -519 -71 -503 -37
rect -445 -71 -429 -37
rect -361 -71 -345 -37
rect -287 -71 -271 -37
rect -203 -71 -187 -37
rect -129 -71 -113 -37
rect -45 -71 -29 -37
rect 29 -71 45 -37
rect 113 -71 129 -37
rect 187 -71 203 -37
rect 271 -71 287 -37
rect 345 -71 361 -37
rect 429 -71 445 -37
rect 503 -71 519 -37
rect 587 -71 603 -37
rect 661 -71 677 -37
rect 745 -71 761 -37
rect -807 -130 -773 -114
rect -807 -1722 -773 -1706
rect -649 -130 -615 -114
rect -649 -1722 -615 -1706
rect -491 -130 -457 -114
rect -491 -1722 -457 -1706
rect -333 -130 -299 -114
rect -333 -1722 -299 -1706
rect -175 -130 -141 -114
rect -175 -1722 -141 -1706
rect -17 -130 17 -114
rect -17 -1722 17 -1706
rect 141 -130 175 -114
rect 141 -1722 175 -1706
rect 299 -130 333 -114
rect 299 -1722 333 -1706
rect 457 -130 491 -114
rect 457 -1722 491 -1706
rect 615 -130 649 -114
rect 615 -1722 649 -1706
rect 773 -130 807 -114
rect 773 -1722 807 -1706
rect -761 -1799 -745 -1765
rect -677 -1799 -661 -1765
rect -603 -1799 -587 -1765
rect -519 -1799 -503 -1765
rect -445 -1799 -429 -1765
rect -361 -1799 -345 -1765
rect -287 -1799 -271 -1765
rect -203 -1799 -187 -1765
rect -129 -1799 -113 -1765
rect -45 -1799 -29 -1765
rect 29 -1799 45 -1765
rect 113 -1799 129 -1765
rect 187 -1799 203 -1765
rect 271 -1799 287 -1765
rect 345 -1799 361 -1765
rect 429 -1799 445 -1765
rect 503 -1799 519 -1765
rect 587 -1799 603 -1765
rect 661 -1799 677 -1765
rect 745 -1799 761 -1765
rect 887 -1867 921 1867
rect -921 -1901 -825 -1867
rect 825 -1901 921 -1867
<< viali >>
rect -745 1765 -677 1799
rect -587 1765 -519 1799
rect -429 1765 -361 1799
rect -271 1765 -203 1799
rect -113 1765 -45 1799
rect 45 1765 113 1799
rect 203 1765 271 1799
rect 361 1765 429 1799
rect 519 1765 587 1799
rect 677 1765 745 1799
rect -807 130 -773 1706
rect -649 130 -615 1706
rect -491 130 -457 1706
rect -333 130 -299 1706
rect -175 130 -141 1706
rect -17 130 17 1706
rect 141 130 175 1706
rect 299 130 333 1706
rect 457 130 491 1706
rect 615 130 649 1706
rect 773 130 807 1706
rect -745 37 -677 71
rect -587 37 -519 71
rect -429 37 -361 71
rect -271 37 -203 71
rect -113 37 -45 71
rect 45 37 113 71
rect 203 37 271 71
rect 361 37 429 71
rect 519 37 587 71
rect 677 37 745 71
rect -745 -71 -677 -37
rect -587 -71 -519 -37
rect -429 -71 -361 -37
rect -271 -71 -203 -37
rect -113 -71 -45 -37
rect 45 -71 113 -37
rect 203 -71 271 -37
rect 361 -71 429 -37
rect 519 -71 587 -37
rect 677 -71 745 -37
rect -807 -1706 -773 -130
rect -649 -1706 -615 -130
rect -491 -1706 -457 -130
rect -333 -1706 -299 -130
rect -175 -1706 -141 -130
rect -17 -1706 17 -130
rect 141 -1706 175 -130
rect 299 -1706 333 -130
rect 457 -1706 491 -130
rect 615 -1706 649 -130
rect 773 -1706 807 -130
rect -745 -1799 -677 -1765
rect -587 -1799 -519 -1765
rect -429 -1799 -361 -1765
rect -271 -1799 -203 -1765
rect -113 -1799 -45 -1765
rect 45 -1799 113 -1765
rect 203 -1799 271 -1765
rect 361 -1799 429 -1765
rect 519 -1799 587 -1765
rect 677 -1799 745 -1765
<< metal1 >>
rect -757 1799 -665 1805
rect -757 1765 -745 1799
rect -677 1765 -665 1799
rect -757 1759 -665 1765
rect -599 1799 -507 1805
rect -599 1765 -587 1799
rect -519 1765 -507 1799
rect -599 1759 -507 1765
rect -441 1799 -349 1805
rect -441 1765 -429 1799
rect -361 1765 -349 1799
rect -441 1759 -349 1765
rect -283 1799 -191 1805
rect -283 1765 -271 1799
rect -203 1765 -191 1799
rect -283 1759 -191 1765
rect -125 1799 -33 1805
rect -125 1765 -113 1799
rect -45 1765 -33 1799
rect -125 1759 -33 1765
rect 33 1799 125 1805
rect 33 1765 45 1799
rect 113 1765 125 1799
rect 33 1759 125 1765
rect 191 1799 283 1805
rect 191 1765 203 1799
rect 271 1765 283 1799
rect 191 1759 283 1765
rect 349 1799 441 1805
rect 349 1765 361 1799
rect 429 1765 441 1799
rect 349 1759 441 1765
rect 507 1799 599 1805
rect 507 1765 519 1799
rect 587 1765 599 1799
rect 507 1759 599 1765
rect 665 1799 757 1805
rect 665 1765 677 1799
rect 745 1765 757 1799
rect 665 1759 757 1765
rect -813 1706 -767 1718
rect -813 130 -807 1706
rect -773 130 -767 1706
rect -813 118 -767 130
rect -655 1706 -609 1718
rect -655 130 -649 1706
rect -615 130 -609 1706
rect -655 118 -609 130
rect -497 1706 -451 1718
rect -497 130 -491 1706
rect -457 130 -451 1706
rect -497 118 -451 130
rect -339 1706 -293 1718
rect -339 130 -333 1706
rect -299 130 -293 1706
rect -339 118 -293 130
rect -181 1706 -135 1718
rect -181 130 -175 1706
rect -141 130 -135 1706
rect -181 118 -135 130
rect -23 1706 23 1718
rect -23 130 -17 1706
rect 17 130 23 1706
rect -23 118 23 130
rect 135 1706 181 1718
rect 135 130 141 1706
rect 175 130 181 1706
rect 135 118 181 130
rect 293 1706 339 1718
rect 293 130 299 1706
rect 333 130 339 1706
rect 293 118 339 130
rect 451 1706 497 1718
rect 451 130 457 1706
rect 491 130 497 1706
rect 451 118 497 130
rect 609 1706 655 1718
rect 609 130 615 1706
rect 649 130 655 1706
rect 609 118 655 130
rect 767 1706 813 1718
rect 767 130 773 1706
rect 807 130 813 1706
rect 767 118 813 130
rect -757 71 -665 77
rect -757 37 -745 71
rect -677 37 -665 71
rect -757 31 -665 37
rect -599 71 -507 77
rect -599 37 -587 71
rect -519 37 -507 71
rect -599 31 -507 37
rect -441 71 -349 77
rect -441 37 -429 71
rect -361 37 -349 71
rect -441 31 -349 37
rect -283 71 -191 77
rect -283 37 -271 71
rect -203 37 -191 71
rect -283 31 -191 37
rect -125 71 -33 77
rect -125 37 -113 71
rect -45 37 -33 71
rect -125 31 -33 37
rect 33 71 125 77
rect 33 37 45 71
rect 113 37 125 71
rect 33 31 125 37
rect 191 71 283 77
rect 191 37 203 71
rect 271 37 283 71
rect 191 31 283 37
rect 349 71 441 77
rect 349 37 361 71
rect 429 37 441 71
rect 349 31 441 37
rect 507 71 599 77
rect 507 37 519 71
rect 587 37 599 71
rect 507 31 599 37
rect 665 71 757 77
rect 665 37 677 71
rect 745 37 757 71
rect 665 31 757 37
rect -757 -37 -665 -31
rect -757 -71 -745 -37
rect -677 -71 -665 -37
rect -757 -77 -665 -71
rect -599 -37 -507 -31
rect -599 -71 -587 -37
rect -519 -71 -507 -37
rect -599 -77 -507 -71
rect -441 -37 -349 -31
rect -441 -71 -429 -37
rect -361 -71 -349 -37
rect -441 -77 -349 -71
rect -283 -37 -191 -31
rect -283 -71 -271 -37
rect -203 -71 -191 -37
rect -283 -77 -191 -71
rect -125 -37 -33 -31
rect -125 -71 -113 -37
rect -45 -71 -33 -37
rect -125 -77 -33 -71
rect 33 -37 125 -31
rect 33 -71 45 -37
rect 113 -71 125 -37
rect 33 -77 125 -71
rect 191 -37 283 -31
rect 191 -71 203 -37
rect 271 -71 283 -37
rect 191 -77 283 -71
rect 349 -37 441 -31
rect 349 -71 361 -37
rect 429 -71 441 -37
rect 349 -77 441 -71
rect 507 -37 599 -31
rect 507 -71 519 -37
rect 587 -71 599 -37
rect 507 -77 599 -71
rect 665 -37 757 -31
rect 665 -71 677 -37
rect 745 -71 757 -37
rect 665 -77 757 -71
rect -813 -130 -767 -118
rect -813 -1706 -807 -130
rect -773 -1706 -767 -130
rect -813 -1718 -767 -1706
rect -655 -130 -609 -118
rect -655 -1706 -649 -130
rect -615 -1706 -609 -130
rect -655 -1718 -609 -1706
rect -497 -130 -451 -118
rect -497 -1706 -491 -130
rect -457 -1706 -451 -130
rect -497 -1718 -451 -1706
rect -339 -130 -293 -118
rect -339 -1706 -333 -130
rect -299 -1706 -293 -130
rect -339 -1718 -293 -1706
rect -181 -130 -135 -118
rect -181 -1706 -175 -130
rect -141 -1706 -135 -130
rect -181 -1718 -135 -1706
rect -23 -130 23 -118
rect -23 -1706 -17 -130
rect 17 -1706 23 -130
rect -23 -1718 23 -1706
rect 135 -130 181 -118
rect 135 -1706 141 -130
rect 175 -1706 181 -130
rect 135 -1718 181 -1706
rect 293 -130 339 -118
rect 293 -1706 299 -130
rect 333 -1706 339 -130
rect 293 -1718 339 -1706
rect 451 -130 497 -118
rect 451 -1706 457 -130
rect 491 -1706 497 -130
rect 451 -1718 497 -1706
rect 609 -130 655 -118
rect 609 -1706 615 -130
rect 649 -1706 655 -130
rect 609 -1718 655 -1706
rect 767 -130 813 -118
rect 767 -1706 773 -130
rect 807 -1706 813 -130
rect 767 -1718 813 -1706
rect -757 -1765 -665 -1759
rect -757 -1799 -745 -1765
rect -677 -1799 -665 -1765
rect -757 -1805 -665 -1799
rect -599 -1765 -507 -1759
rect -599 -1799 -587 -1765
rect -519 -1799 -507 -1765
rect -599 -1805 -507 -1799
rect -441 -1765 -349 -1759
rect -441 -1799 -429 -1765
rect -361 -1799 -349 -1765
rect -441 -1805 -349 -1799
rect -283 -1765 -191 -1759
rect -283 -1799 -271 -1765
rect -203 -1799 -191 -1765
rect -283 -1805 -191 -1799
rect -125 -1765 -33 -1759
rect -125 -1799 -113 -1765
rect -45 -1799 -33 -1765
rect -125 -1805 -33 -1799
rect 33 -1765 125 -1759
rect 33 -1799 45 -1765
rect 113 -1799 125 -1765
rect 33 -1805 125 -1799
rect 191 -1765 283 -1759
rect 191 -1799 203 -1765
rect 271 -1799 283 -1765
rect 191 -1805 283 -1799
rect 349 -1765 441 -1759
rect 349 -1799 361 -1765
rect 429 -1799 441 -1765
rect 349 -1805 441 -1799
rect 507 -1765 599 -1759
rect 507 -1799 519 -1765
rect 587 -1799 599 -1765
rect 507 -1805 599 -1799
rect 665 -1765 757 -1759
rect 665 -1799 677 -1765
rect 745 -1799 757 -1765
rect 665 -1805 757 -1799
<< properties >>
string FIXED_BBOX -904 -1884 904 1884
string gencell sky130_fd_pr__pfet_01v8_lvt
string library sky130
string parameters w 8 l 0.5 m 2 nf 10 diffcov 100 polycov 100 guard 1 glc 0 grc 0 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.35 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
