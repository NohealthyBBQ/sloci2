magic
tech sky130A
magscale 1 2
timestamp 1671745787
<< error_p >>
rect -461 1217 -403 1223
rect -269 1217 -211 1223
rect -77 1217 -19 1223
rect 115 1217 173 1223
rect 307 1217 365 1223
rect -461 1183 -449 1217
rect -269 1183 -257 1217
rect -77 1183 -65 1217
rect 115 1183 127 1217
rect 307 1183 319 1217
rect -461 1177 -403 1183
rect -269 1177 -211 1183
rect -77 1177 -19 1183
rect 115 1177 173 1183
rect 307 1177 365 1183
rect -365 907 -307 913
rect -173 907 -115 913
rect 19 907 77 913
rect 211 907 269 913
rect 403 907 461 913
rect -365 873 -353 907
rect -173 873 -161 907
rect 19 873 31 907
rect 211 873 223 907
rect 403 873 415 907
rect -365 867 -307 873
rect -173 867 -115 873
rect 19 867 77 873
rect 211 867 269 873
rect 403 867 461 873
rect -365 799 -307 805
rect -173 799 -115 805
rect 19 799 77 805
rect 211 799 269 805
rect 403 799 461 805
rect -365 765 -353 799
rect -173 765 -161 799
rect 19 765 31 799
rect 211 765 223 799
rect 403 765 415 799
rect -365 759 -307 765
rect -173 759 -115 765
rect 19 759 77 765
rect 211 759 269 765
rect 403 759 461 765
rect -461 489 -403 495
rect -269 489 -211 495
rect -77 489 -19 495
rect 115 489 173 495
rect 307 489 365 495
rect -461 455 -449 489
rect -269 455 -257 489
rect -77 455 -65 489
rect 115 455 127 489
rect 307 455 319 489
rect -461 449 -403 455
rect -269 449 -211 455
rect -77 449 -19 455
rect 115 449 173 455
rect 307 449 365 455
rect -461 381 -403 387
rect -269 381 -211 387
rect -77 381 -19 387
rect 115 381 173 387
rect 307 381 365 387
rect -461 347 -449 381
rect -269 347 -257 381
rect -77 347 -65 381
rect 115 347 127 381
rect 307 347 319 381
rect -461 341 -403 347
rect -269 341 -211 347
rect -77 341 -19 347
rect 115 341 173 347
rect 307 341 365 347
rect -365 71 -307 77
rect -173 71 -115 77
rect 19 71 77 77
rect 211 71 269 77
rect 403 71 461 77
rect -365 37 -353 71
rect -173 37 -161 71
rect 19 37 31 71
rect 211 37 223 71
rect 403 37 415 71
rect -365 31 -307 37
rect -173 31 -115 37
rect 19 31 77 37
rect 211 31 269 37
rect 403 31 461 37
rect -365 -37 -307 -31
rect -173 -37 -115 -31
rect 19 -37 77 -31
rect 211 -37 269 -31
rect 403 -37 461 -31
rect -365 -71 -353 -37
rect -173 -71 -161 -37
rect 19 -71 31 -37
rect 211 -71 223 -37
rect 403 -71 415 -37
rect -365 -77 -307 -71
rect -173 -77 -115 -71
rect 19 -77 77 -71
rect 211 -77 269 -71
rect 403 -77 461 -71
rect -461 -347 -403 -341
rect -269 -347 -211 -341
rect -77 -347 -19 -341
rect 115 -347 173 -341
rect 307 -347 365 -341
rect -461 -381 -449 -347
rect -269 -381 -257 -347
rect -77 -381 -65 -347
rect 115 -381 127 -347
rect 307 -381 319 -347
rect -461 -387 -403 -381
rect -269 -387 -211 -381
rect -77 -387 -19 -381
rect 115 -387 173 -381
rect 307 -387 365 -381
rect -461 -455 -403 -449
rect -269 -455 -211 -449
rect -77 -455 -19 -449
rect 115 -455 173 -449
rect 307 -455 365 -449
rect -461 -489 -449 -455
rect -269 -489 -257 -455
rect -77 -489 -65 -455
rect 115 -489 127 -455
rect 307 -489 319 -455
rect -461 -495 -403 -489
rect -269 -495 -211 -489
rect -77 -495 -19 -489
rect 115 -495 173 -489
rect 307 -495 365 -489
rect -365 -765 -307 -759
rect -173 -765 -115 -759
rect 19 -765 77 -759
rect 211 -765 269 -759
rect 403 -765 461 -759
rect -365 -799 -353 -765
rect -173 -799 -161 -765
rect 19 -799 31 -765
rect 211 -799 223 -765
rect 403 -799 415 -765
rect -365 -805 -307 -799
rect -173 -805 -115 -799
rect 19 -805 77 -799
rect 211 -805 269 -799
rect 403 -805 461 -799
rect -365 -873 -307 -867
rect -173 -873 -115 -867
rect 19 -873 77 -867
rect 211 -873 269 -867
rect 403 -873 461 -867
rect -365 -907 -353 -873
rect -173 -907 -161 -873
rect 19 -907 31 -873
rect 211 -907 223 -873
rect 403 -907 415 -873
rect -365 -913 -307 -907
rect -173 -913 -115 -907
rect 19 -913 77 -907
rect 211 -913 269 -907
rect 403 -913 461 -907
rect -461 -1183 -403 -1177
rect -269 -1183 -211 -1177
rect -77 -1183 -19 -1177
rect 115 -1183 173 -1177
rect 307 -1183 365 -1177
rect -461 -1217 -449 -1183
rect -269 -1217 -257 -1183
rect -77 -1217 -65 -1183
rect 115 -1217 127 -1183
rect 307 -1217 319 -1183
rect -461 -1223 -403 -1217
rect -269 -1223 -211 -1217
rect -77 -1223 -19 -1217
rect 115 -1223 173 -1217
rect 307 -1223 365 -1217
<< pwell >>
rect -647 -1355 647 1355
<< nmoslvt >>
rect -447 945 -417 1145
rect -351 945 -321 1145
rect -255 945 -225 1145
rect -159 945 -129 1145
rect -63 945 -33 1145
rect 33 945 63 1145
rect 129 945 159 1145
rect 225 945 255 1145
rect 321 945 351 1145
rect 417 945 447 1145
rect -447 527 -417 727
rect -351 527 -321 727
rect -255 527 -225 727
rect -159 527 -129 727
rect -63 527 -33 727
rect 33 527 63 727
rect 129 527 159 727
rect 225 527 255 727
rect 321 527 351 727
rect 417 527 447 727
rect -447 109 -417 309
rect -351 109 -321 309
rect -255 109 -225 309
rect -159 109 -129 309
rect -63 109 -33 309
rect 33 109 63 309
rect 129 109 159 309
rect 225 109 255 309
rect 321 109 351 309
rect 417 109 447 309
rect -447 -309 -417 -109
rect -351 -309 -321 -109
rect -255 -309 -225 -109
rect -159 -309 -129 -109
rect -63 -309 -33 -109
rect 33 -309 63 -109
rect 129 -309 159 -109
rect 225 -309 255 -109
rect 321 -309 351 -109
rect 417 -309 447 -109
rect -447 -727 -417 -527
rect -351 -727 -321 -527
rect -255 -727 -225 -527
rect -159 -727 -129 -527
rect -63 -727 -33 -527
rect 33 -727 63 -527
rect 129 -727 159 -527
rect 225 -727 255 -527
rect 321 -727 351 -527
rect 417 -727 447 -527
rect -447 -1145 -417 -945
rect -351 -1145 -321 -945
rect -255 -1145 -225 -945
rect -159 -1145 -129 -945
rect -63 -1145 -33 -945
rect 33 -1145 63 -945
rect 129 -1145 159 -945
rect 225 -1145 255 -945
rect 321 -1145 351 -945
rect 417 -1145 447 -945
<< ndiff >>
rect -509 1133 -447 1145
rect -509 957 -497 1133
rect -463 957 -447 1133
rect -509 945 -447 957
rect -417 1133 -351 1145
rect -417 957 -401 1133
rect -367 957 -351 1133
rect -417 945 -351 957
rect -321 1133 -255 1145
rect -321 957 -305 1133
rect -271 957 -255 1133
rect -321 945 -255 957
rect -225 1133 -159 1145
rect -225 957 -209 1133
rect -175 957 -159 1133
rect -225 945 -159 957
rect -129 1133 -63 1145
rect -129 957 -113 1133
rect -79 957 -63 1133
rect -129 945 -63 957
rect -33 1133 33 1145
rect -33 957 -17 1133
rect 17 957 33 1133
rect -33 945 33 957
rect 63 1133 129 1145
rect 63 957 79 1133
rect 113 957 129 1133
rect 63 945 129 957
rect 159 1133 225 1145
rect 159 957 175 1133
rect 209 957 225 1133
rect 159 945 225 957
rect 255 1133 321 1145
rect 255 957 271 1133
rect 305 957 321 1133
rect 255 945 321 957
rect 351 1133 417 1145
rect 351 957 367 1133
rect 401 957 417 1133
rect 351 945 417 957
rect 447 1133 509 1145
rect 447 957 463 1133
rect 497 957 509 1133
rect 447 945 509 957
rect -509 715 -447 727
rect -509 539 -497 715
rect -463 539 -447 715
rect -509 527 -447 539
rect -417 715 -351 727
rect -417 539 -401 715
rect -367 539 -351 715
rect -417 527 -351 539
rect -321 715 -255 727
rect -321 539 -305 715
rect -271 539 -255 715
rect -321 527 -255 539
rect -225 715 -159 727
rect -225 539 -209 715
rect -175 539 -159 715
rect -225 527 -159 539
rect -129 715 -63 727
rect -129 539 -113 715
rect -79 539 -63 715
rect -129 527 -63 539
rect -33 715 33 727
rect -33 539 -17 715
rect 17 539 33 715
rect -33 527 33 539
rect 63 715 129 727
rect 63 539 79 715
rect 113 539 129 715
rect 63 527 129 539
rect 159 715 225 727
rect 159 539 175 715
rect 209 539 225 715
rect 159 527 225 539
rect 255 715 321 727
rect 255 539 271 715
rect 305 539 321 715
rect 255 527 321 539
rect 351 715 417 727
rect 351 539 367 715
rect 401 539 417 715
rect 351 527 417 539
rect 447 715 509 727
rect 447 539 463 715
rect 497 539 509 715
rect 447 527 509 539
rect -509 297 -447 309
rect -509 121 -497 297
rect -463 121 -447 297
rect -509 109 -447 121
rect -417 297 -351 309
rect -417 121 -401 297
rect -367 121 -351 297
rect -417 109 -351 121
rect -321 297 -255 309
rect -321 121 -305 297
rect -271 121 -255 297
rect -321 109 -255 121
rect -225 297 -159 309
rect -225 121 -209 297
rect -175 121 -159 297
rect -225 109 -159 121
rect -129 297 -63 309
rect -129 121 -113 297
rect -79 121 -63 297
rect -129 109 -63 121
rect -33 297 33 309
rect -33 121 -17 297
rect 17 121 33 297
rect -33 109 33 121
rect 63 297 129 309
rect 63 121 79 297
rect 113 121 129 297
rect 63 109 129 121
rect 159 297 225 309
rect 159 121 175 297
rect 209 121 225 297
rect 159 109 225 121
rect 255 297 321 309
rect 255 121 271 297
rect 305 121 321 297
rect 255 109 321 121
rect 351 297 417 309
rect 351 121 367 297
rect 401 121 417 297
rect 351 109 417 121
rect 447 297 509 309
rect 447 121 463 297
rect 497 121 509 297
rect 447 109 509 121
rect -509 -121 -447 -109
rect -509 -297 -497 -121
rect -463 -297 -447 -121
rect -509 -309 -447 -297
rect -417 -121 -351 -109
rect -417 -297 -401 -121
rect -367 -297 -351 -121
rect -417 -309 -351 -297
rect -321 -121 -255 -109
rect -321 -297 -305 -121
rect -271 -297 -255 -121
rect -321 -309 -255 -297
rect -225 -121 -159 -109
rect -225 -297 -209 -121
rect -175 -297 -159 -121
rect -225 -309 -159 -297
rect -129 -121 -63 -109
rect -129 -297 -113 -121
rect -79 -297 -63 -121
rect -129 -309 -63 -297
rect -33 -121 33 -109
rect -33 -297 -17 -121
rect 17 -297 33 -121
rect -33 -309 33 -297
rect 63 -121 129 -109
rect 63 -297 79 -121
rect 113 -297 129 -121
rect 63 -309 129 -297
rect 159 -121 225 -109
rect 159 -297 175 -121
rect 209 -297 225 -121
rect 159 -309 225 -297
rect 255 -121 321 -109
rect 255 -297 271 -121
rect 305 -297 321 -121
rect 255 -309 321 -297
rect 351 -121 417 -109
rect 351 -297 367 -121
rect 401 -297 417 -121
rect 351 -309 417 -297
rect 447 -121 509 -109
rect 447 -297 463 -121
rect 497 -297 509 -121
rect 447 -309 509 -297
rect -509 -539 -447 -527
rect -509 -715 -497 -539
rect -463 -715 -447 -539
rect -509 -727 -447 -715
rect -417 -539 -351 -527
rect -417 -715 -401 -539
rect -367 -715 -351 -539
rect -417 -727 -351 -715
rect -321 -539 -255 -527
rect -321 -715 -305 -539
rect -271 -715 -255 -539
rect -321 -727 -255 -715
rect -225 -539 -159 -527
rect -225 -715 -209 -539
rect -175 -715 -159 -539
rect -225 -727 -159 -715
rect -129 -539 -63 -527
rect -129 -715 -113 -539
rect -79 -715 -63 -539
rect -129 -727 -63 -715
rect -33 -539 33 -527
rect -33 -715 -17 -539
rect 17 -715 33 -539
rect -33 -727 33 -715
rect 63 -539 129 -527
rect 63 -715 79 -539
rect 113 -715 129 -539
rect 63 -727 129 -715
rect 159 -539 225 -527
rect 159 -715 175 -539
rect 209 -715 225 -539
rect 159 -727 225 -715
rect 255 -539 321 -527
rect 255 -715 271 -539
rect 305 -715 321 -539
rect 255 -727 321 -715
rect 351 -539 417 -527
rect 351 -715 367 -539
rect 401 -715 417 -539
rect 351 -727 417 -715
rect 447 -539 509 -527
rect 447 -715 463 -539
rect 497 -715 509 -539
rect 447 -727 509 -715
rect -509 -957 -447 -945
rect -509 -1133 -497 -957
rect -463 -1133 -447 -957
rect -509 -1145 -447 -1133
rect -417 -957 -351 -945
rect -417 -1133 -401 -957
rect -367 -1133 -351 -957
rect -417 -1145 -351 -1133
rect -321 -957 -255 -945
rect -321 -1133 -305 -957
rect -271 -1133 -255 -957
rect -321 -1145 -255 -1133
rect -225 -957 -159 -945
rect -225 -1133 -209 -957
rect -175 -1133 -159 -957
rect -225 -1145 -159 -1133
rect -129 -957 -63 -945
rect -129 -1133 -113 -957
rect -79 -1133 -63 -957
rect -129 -1145 -63 -1133
rect -33 -957 33 -945
rect -33 -1133 -17 -957
rect 17 -1133 33 -957
rect -33 -1145 33 -1133
rect 63 -957 129 -945
rect 63 -1133 79 -957
rect 113 -1133 129 -957
rect 63 -1145 129 -1133
rect 159 -957 225 -945
rect 159 -1133 175 -957
rect 209 -1133 225 -957
rect 159 -1145 225 -1133
rect 255 -957 321 -945
rect 255 -1133 271 -957
rect 305 -1133 321 -957
rect 255 -1145 321 -1133
rect 351 -957 417 -945
rect 351 -1133 367 -957
rect 401 -1133 417 -957
rect 351 -1145 417 -1133
rect 447 -957 509 -945
rect 447 -1133 463 -957
rect 497 -1133 509 -957
rect 447 -1145 509 -1133
<< ndiffc >>
rect -497 957 -463 1133
rect -401 957 -367 1133
rect -305 957 -271 1133
rect -209 957 -175 1133
rect -113 957 -79 1133
rect -17 957 17 1133
rect 79 957 113 1133
rect 175 957 209 1133
rect 271 957 305 1133
rect 367 957 401 1133
rect 463 957 497 1133
rect -497 539 -463 715
rect -401 539 -367 715
rect -305 539 -271 715
rect -209 539 -175 715
rect -113 539 -79 715
rect -17 539 17 715
rect 79 539 113 715
rect 175 539 209 715
rect 271 539 305 715
rect 367 539 401 715
rect 463 539 497 715
rect -497 121 -463 297
rect -401 121 -367 297
rect -305 121 -271 297
rect -209 121 -175 297
rect -113 121 -79 297
rect -17 121 17 297
rect 79 121 113 297
rect 175 121 209 297
rect 271 121 305 297
rect 367 121 401 297
rect 463 121 497 297
rect -497 -297 -463 -121
rect -401 -297 -367 -121
rect -305 -297 -271 -121
rect -209 -297 -175 -121
rect -113 -297 -79 -121
rect -17 -297 17 -121
rect 79 -297 113 -121
rect 175 -297 209 -121
rect 271 -297 305 -121
rect 367 -297 401 -121
rect 463 -297 497 -121
rect -497 -715 -463 -539
rect -401 -715 -367 -539
rect -305 -715 -271 -539
rect -209 -715 -175 -539
rect -113 -715 -79 -539
rect -17 -715 17 -539
rect 79 -715 113 -539
rect 175 -715 209 -539
rect 271 -715 305 -539
rect 367 -715 401 -539
rect 463 -715 497 -539
rect -497 -1133 -463 -957
rect -401 -1133 -367 -957
rect -305 -1133 -271 -957
rect -209 -1133 -175 -957
rect -113 -1133 -79 -957
rect -17 -1133 17 -957
rect 79 -1133 113 -957
rect 175 -1133 209 -957
rect 271 -1133 305 -957
rect 367 -1133 401 -957
rect 463 -1133 497 -957
<< psubdiff >>
rect -611 1285 -515 1319
rect 515 1285 611 1319
rect -611 1223 -577 1285
rect 577 1223 611 1285
rect -611 -1285 -577 -1223
rect 577 -1285 611 -1223
rect -611 -1319 -515 -1285
rect 515 -1319 611 -1285
<< psubdiffcont >>
rect -515 1285 515 1319
rect -611 -1223 -577 1223
rect 577 -1223 611 1223
rect -515 -1319 515 -1285
<< poly >>
rect -465 1217 -399 1233
rect -465 1183 -449 1217
rect -415 1183 -399 1217
rect -465 1167 -399 1183
rect -273 1217 -207 1233
rect -273 1183 -257 1217
rect -223 1183 -207 1217
rect -447 1145 -417 1167
rect -351 1145 -321 1171
rect -273 1167 -207 1183
rect -81 1217 -15 1233
rect -81 1183 -65 1217
rect -31 1183 -15 1217
rect -255 1145 -225 1167
rect -159 1145 -129 1171
rect -81 1167 -15 1183
rect 111 1217 177 1233
rect 111 1183 127 1217
rect 161 1183 177 1217
rect -63 1145 -33 1167
rect 33 1145 63 1171
rect 111 1167 177 1183
rect 303 1217 369 1233
rect 303 1183 319 1217
rect 353 1183 369 1217
rect 129 1145 159 1167
rect 225 1145 255 1171
rect 303 1167 369 1183
rect 321 1145 351 1167
rect 417 1145 447 1171
rect -447 919 -417 945
rect -351 923 -321 945
rect -369 907 -303 923
rect -255 919 -225 945
rect -159 923 -129 945
rect -369 873 -353 907
rect -319 873 -303 907
rect -369 857 -303 873
rect -177 907 -111 923
rect -63 919 -33 945
rect 33 923 63 945
rect -177 873 -161 907
rect -127 873 -111 907
rect -177 857 -111 873
rect 15 907 81 923
rect 129 919 159 945
rect 225 923 255 945
rect 15 873 31 907
rect 65 873 81 907
rect 15 857 81 873
rect 207 907 273 923
rect 321 919 351 945
rect 417 923 447 945
rect 207 873 223 907
rect 257 873 273 907
rect 207 857 273 873
rect 399 907 465 923
rect 399 873 415 907
rect 449 873 465 907
rect 399 857 465 873
rect -369 799 -303 815
rect -369 765 -353 799
rect -319 765 -303 799
rect -447 727 -417 753
rect -369 749 -303 765
rect -177 799 -111 815
rect -177 765 -161 799
rect -127 765 -111 799
rect -351 727 -321 749
rect -255 727 -225 753
rect -177 749 -111 765
rect 15 799 81 815
rect 15 765 31 799
rect 65 765 81 799
rect -159 727 -129 749
rect -63 727 -33 753
rect 15 749 81 765
rect 207 799 273 815
rect 207 765 223 799
rect 257 765 273 799
rect 33 727 63 749
rect 129 727 159 753
rect 207 749 273 765
rect 399 799 465 815
rect 399 765 415 799
rect 449 765 465 799
rect 225 727 255 749
rect 321 727 351 753
rect 399 749 465 765
rect 417 727 447 749
rect -447 505 -417 527
rect -465 489 -399 505
rect -351 501 -321 527
rect -255 505 -225 527
rect -465 455 -449 489
rect -415 455 -399 489
rect -465 439 -399 455
rect -273 489 -207 505
rect -159 501 -129 527
rect -63 505 -33 527
rect -273 455 -257 489
rect -223 455 -207 489
rect -273 439 -207 455
rect -81 489 -15 505
rect 33 501 63 527
rect 129 505 159 527
rect -81 455 -65 489
rect -31 455 -15 489
rect -81 439 -15 455
rect 111 489 177 505
rect 225 501 255 527
rect 321 505 351 527
rect 111 455 127 489
rect 161 455 177 489
rect 111 439 177 455
rect 303 489 369 505
rect 417 501 447 527
rect 303 455 319 489
rect 353 455 369 489
rect 303 439 369 455
rect -465 381 -399 397
rect -465 347 -449 381
rect -415 347 -399 381
rect -465 331 -399 347
rect -273 381 -207 397
rect -273 347 -257 381
rect -223 347 -207 381
rect -447 309 -417 331
rect -351 309 -321 335
rect -273 331 -207 347
rect -81 381 -15 397
rect -81 347 -65 381
rect -31 347 -15 381
rect -255 309 -225 331
rect -159 309 -129 335
rect -81 331 -15 347
rect 111 381 177 397
rect 111 347 127 381
rect 161 347 177 381
rect -63 309 -33 331
rect 33 309 63 335
rect 111 331 177 347
rect 303 381 369 397
rect 303 347 319 381
rect 353 347 369 381
rect 129 309 159 331
rect 225 309 255 335
rect 303 331 369 347
rect 321 309 351 331
rect 417 309 447 335
rect -447 83 -417 109
rect -351 87 -321 109
rect -369 71 -303 87
rect -255 83 -225 109
rect -159 87 -129 109
rect -369 37 -353 71
rect -319 37 -303 71
rect -369 21 -303 37
rect -177 71 -111 87
rect -63 83 -33 109
rect 33 87 63 109
rect -177 37 -161 71
rect -127 37 -111 71
rect -177 21 -111 37
rect 15 71 81 87
rect 129 83 159 109
rect 225 87 255 109
rect 15 37 31 71
rect 65 37 81 71
rect 15 21 81 37
rect 207 71 273 87
rect 321 83 351 109
rect 417 87 447 109
rect 207 37 223 71
rect 257 37 273 71
rect 207 21 273 37
rect 399 71 465 87
rect 399 37 415 71
rect 449 37 465 71
rect 399 21 465 37
rect -369 -37 -303 -21
rect -369 -71 -353 -37
rect -319 -71 -303 -37
rect -447 -109 -417 -83
rect -369 -87 -303 -71
rect -177 -37 -111 -21
rect -177 -71 -161 -37
rect -127 -71 -111 -37
rect -351 -109 -321 -87
rect -255 -109 -225 -83
rect -177 -87 -111 -71
rect 15 -37 81 -21
rect 15 -71 31 -37
rect 65 -71 81 -37
rect -159 -109 -129 -87
rect -63 -109 -33 -83
rect 15 -87 81 -71
rect 207 -37 273 -21
rect 207 -71 223 -37
rect 257 -71 273 -37
rect 33 -109 63 -87
rect 129 -109 159 -83
rect 207 -87 273 -71
rect 399 -37 465 -21
rect 399 -71 415 -37
rect 449 -71 465 -37
rect 225 -109 255 -87
rect 321 -109 351 -83
rect 399 -87 465 -71
rect 417 -109 447 -87
rect -447 -331 -417 -309
rect -465 -347 -399 -331
rect -351 -335 -321 -309
rect -255 -331 -225 -309
rect -465 -381 -449 -347
rect -415 -381 -399 -347
rect -465 -397 -399 -381
rect -273 -347 -207 -331
rect -159 -335 -129 -309
rect -63 -331 -33 -309
rect -273 -381 -257 -347
rect -223 -381 -207 -347
rect -273 -397 -207 -381
rect -81 -347 -15 -331
rect 33 -335 63 -309
rect 129 -331 159 -309
rect -81 -381 -65 -347
rect -31 -381 -15 -347
rect -81 -397 -15 -381
rect 111 -347 177 -331
rect 225 -335 255 -309
rect 321 -331 351 -309
rect 111 -381 127 -347
rect 161 -381 177 -347
rect 111 -397 177 -381
rect 303 -347 369 -331
rect 417 -335 447 -309
rect 303 -381 319 -347
rect 353 -381 369 -347
rect 303 -397 369 -381
rect -465 -455 -399 -439
rect -465 -489 -449 -455
rect -415 -489 -399 -455
rect -465 -505 -399 -489
rect -273 -455 -207 -439
rect -273 -489 -257 -455
rect -223 -489 -207 -455
rect -447 -527 -417 -505
rect -351 -527 -321 -501
rect -273 -505 -207 -489
rect -81 -455 -15 -439
rect -81 -489 -65 -455
rect -31 -489 -15 -455
rect -255 -527 -225 -505
rect -159 -527 -129 -501
rect -81 -505 -15 -489
rect 111 -455 177 -439
rect 111 -489 127 -455
rect 161 -489 177 -455
rect -63 -527 -33 -505
rect 33 -527 63 -501
rect 111 -505 177 -489
rect 303 -455 369 -439
rect 303 -489 319 -455
rect 353 -489 369 -455
rect 129 -527 159 -505
rect 225 -527 255 -501
rect 303 -505 369 -489
rect 321 -527 351 -505
rect 417 -527 447 -501
rect -447 -753 -417 -727
rect -351 -749 -321 -727
rect -369 -765 -303 -749
rect -255 -753 -225 -727
rect -159 -749 -129 -727
rect -369 -799 -353 -765
rect -319 -799 -303 -765
rect -369 -815 -303 -799
rect -177 -765 -111 -749
rect -63 -753 -33 -727
rect 33 -749 63 -727
rect -177 -799 -161 -765
rect -127 -799 -111 -765
rect -177 -815 -111 -799
rect 15 -765 81 -749
rect 129 -753 159 -727
rect 225 -749 255 -727
rect 15 -799 31 -765
rect 65 -799 81 -765
rect 15 -815 81 -799
rect 207 -765 273 -749
rect 321 -753 351 -727
rect 417 -749 447 -727
rect 207 -799 223 -765
rect 257 -799 273 -765
rect 207 -815 273 -799
rect 399 -765 465 -749
rect 399 -799 415 -765
rect 449 -799 465 -765
rect 399 -815 465 -799
rect -369 -873 -303 -857
rect -369 -907 -353 -873
rect -319 -907 -303 -873
rect -447 -945 -417 -919
rect -369 -923 -303 -907
rect -177 -873 -111 -857
rect -177 -907 -161 -873
rect -127 -907 -111 -873
rect -351 -945 -321 -923
rect -255 -945 -225 -919
rect -177 -923 -111 -907
rect 15 -873 81 -857
rect 15 -907 31 -873
rect 65 -907 81 -873
rect -159 -945 -129 -923
rect -63 -945 -33 -919
rect 15 -923 81 -907
rect 207 -873 273 -857
rect 207 -907 223 -873
rect 257 -907 273 -873
rect 33 -945 63 -923
rect 129 -945 159 -919
rect 207 -923 273 -907
rect 399 -873 465 -857
rect 399 -907 415 -873
rect 449 -907 465 -873
rect 225 -945 255 -923
rect 321 -945 351 -919
rect 399 -923 465 -907
rect 417 -945 447 -923
rect -447 -1167 -417 -1145
rect -465 -1183 -399 -1167
rect -351 -1171 -321 -1145
rect -255 -1167 -225 -1145
rect -465 -1217 -449 -1183
rect -415 -1217 -399 -1183
rect -465 -1233 -399 -1217
rect -273 -1183 -207 -1167
rect -159 -1171 -129 -1145
rect -63 -1167 -33 -1145
rect -273 -1217 -257 -1183
rect -223 -1217 -207 -1183
rect -273 -1233 -207 -1217
rect -81 -1183 -15 -1167
rect 33 -1171 63 -1145
rect 129 -1167 159 -1145
rect -81 -1217 -65 -1183
rect -31 -1217 -15 -1183
rect -81 -1233 -15 -1217
rect 111 -1183 177 -1167
rect 225 -1171 255 -1145
rect 321 -1167 351 -1145
rect 111 -1217 127 -1183
rect 161 -1217 177 -1183
rect 111 -1233 177 -1217
rect 303 -1183 369 -1167
rect 417 -1171 447 -1145
rect 303 -1217 319 -1183
rect 353 -1217 369 -1183
rect 303 -1233 369 -1217
<< polycont >>
rect -449 1183 -415 1217
rect -257 1183 -223 1217
rect -65 1183 -31 1217
rect 127 1183 161 1217
rect 319 1183 353 1217
rect -353 873 -319 907
rect -161 873 -127 907
rect 31 873 65 907
rect 223 873 257 907
rect 415 873 449 907
rect -353 765 -319 799
rect -161 765 -127 799
rect 31 765 65 799
rect 223 765 257 799
rect 415 765 449 799
rect -449 455 -415 489
rect -257 455 -223 489
rect -65 455 -31 489
rect 127 455 161 489
rect 319 455 353 489
rect -449 347 -415 381
rect -257 347 -223 381
rect -65 347 -31 381
rect 127 347 161 381
rect 319 347 353 381
rect -353 37 -319 71
rect -161 37 -127 71
rect 31 37 65 71
rect 223 37 257 71
rect 415 37 449 71
rect -353 -71 -319 -37
rect -161 -71 -127 -37
rect 31 -71 65 -37
rect 223 -71 257 -37
rect 415 -71 449 -37
rect -449 -381 -415 -347
rect -257 -381 -223 -347
rect -65 -381 -31 -347
rect 127 -381 161 -347
rect 319 -381 353 -347
rect -449 -489 -415 -455
rect -257 -489 -223 -455
rect -65 -489 -31 -455
rect 127 -489 161 -455
rect 319 -489 353 -455
rect -353 -799 -319 -765
rect -161 -799 -127 -765
rect 31 -799 65 -765
rect 223 -799 257 -765
rect 415 -799 449 -765
rect -353 -907 -319 -873
rect -161 -907 -127 -873
rect 31 -907 65 -873
rect 223 -907 257 -873
rect 415 -907 449 -873
rect -449 -1217 -415 -1183
rect -257 -1217 -223 -1183
rect -65 -1217 -31 -1183
rect 127 -1217 161 -1183
rect 319 -1217 353 -1183
<< locali >>
rect -611 1285 -515 1319
rect 515 1285 611 1319
rect -611 1223 -577 1285
rect 577 1223 611 1285
rect -465 1183 -449 1217
rect -415 1183 -399 1217
rect -273 1183 -257 1217
rect -223 1183 -207 1217
rect -81 1183 -65 1217
rect -31 1183 -15 1217
rect 111 1183 127 1217
rect 161 1183 177 1217
rect 303 1183 319 1217
rect 353 1183 369 1217
rect -497 1133 -463 1149
rect -497 941 -463 957
rect -401 1133 -367 1149
rect -401 941 -367 957
rect -305 1133 -271 1149
rect -305 941 -271 957
rect -209 1133 -175 1149
rect -209 941 -175 957
rect -113 1133 -79 1149
rect -113 941 -79 957
rect -17 1133 17 1149
rect -17 941 17 957
rect 79 1133 113 1149
rect 79 941 113 957
rect 175 1133 209 1149
rect 175 941 209 957
rect 271 1133 305 1149
rect 271 941 305 957
rect 367 1133 401 1149
rect 367 941 401 957
rect 463 1133 497 1149
rect 463 941 497 957
rect -369 873 -353 907
rect -319 873 -303 907
rect -177 873 -161 907
rect -127 873 -111 907
rect 15 873 31 907
rect 65 873 81 907
rect 207 873 223 907
rect 257 873 273 907
rect 399 873 415 907
rect 449 873 465 907
rect -369 765 -353 799
rect -319 765 -303 799
rect -177 765 -161 799
rect -127 765 -111 799
rect 15 765 31 799
rect 65 765 81 799
rect 207 765 223 799
rect 257 765 273 799
rect 399 765 415 799
rect 449 765 465 799
rect -497 715 -463 731
rect -497 523 -463 539
rect -401 715 -367 731
rect -401 523 -367 539
rect -305 715 -271 731
rect -305 523 -271 539
rect -209 715 -175 731
rect -209 523 -175 539
rect -113 715 -79 731
rect -113 523 -79 539
rect -17 715 17 731
rect -17 523 17 539
rect 79 715 113 731
rect 79 523 113 539
rect 175 715 209 731
rect 175 523 209 539
rect 271 715 305 731
rect 271 523 305 539
rect 367 715 401 731
rect 367 523 401 539
rect 463 715 497 731
rect 463 523 497 539
rect -465 455 -449 489
rect -415 455 -399 489
rect -273 455 -257 489
rect -223 455 -207 489
rect -81 455 -65 489
rect -31 455 -15 489
rect 111 455 127 489
rect 161 455 177 489
rect 303 455 319 489
rect 353 455 369 489
rect -465 347 -449 381
rect -415 347 -399 381
rect -273 347 -257 381
rect -223 347 -207 381
rect -81 347 -65 381
rect -31 347 -15 381
rect 111 347 127 381
rect 161 347 177 381
rect 303 347 319 381
rect 353 347 369 381
rect -497 297 -463 313
rect -497 105 -463 121
rect -401 297 -367 313
rect -401 105 -367 121
rect -305 297 -271 313
rect -305 105 -271 121
rect -209 297 -175 313
rect -209 105 -175 121
rect -113 297 -79 313
rect -113 105 -79 121
rect -17 297 17 313
rect -17 105 17 121
rect 79 297 113 313
rect 79 105 113 121
rect 175 297 209 313
rect 175 105 209 121
rect 271 297 305 313
rect 271 105 305 121
rect 367 297 401 313
rect 367 105 401 121
rect 463 297 497 313
rect 463 105 497 121
rect -369 37 -353 71
rect -319 37 -303 71
rect -177 37 -161 71
rect -127 37 -111 71
rect 15 37 31 71
rect 65 37 81 71
rect 207 37 223 71
rect 257 37 273 71
rect 399 37 415 71
rect 449 37 465 71
rect -369 -71 -353 -37
rect -319 -71 -303 -37
rect -177 -71 -161 -37
rect -127 -71 -111 -37
rect 15 -71 31 -37
rect 65 -71 81 -37
rect 207 -71 223 -37
rect 257 -71 273 -37
rect 399 -71 415 -37
rect 449 -71 465 -37
rect -497 -121 -463 -105
rect -497 -313 -463 -297
rect -401 -121 -367 -105
rect -401 -313 -367 -297
rect -305 -121 -271 -105
rect -305 -313 -271 -297
rect -209 -121 -175 -105
rect -209 -313 -175 -297
rect -113 -121 -79 -105
rect -113 -313 -79 -297
rect -17 -121 17 -105
rect -17 -313 17 -297
rect 79 -121 113 -105
rect 79 -313 113 -297
rect 175 -121 209 -105
rect 175 -313 209 -297
rect 271 -121 305 -105
rect 271 -313 305 -297
rect 367 -121 401 -105
rect 367 -313 401 -297
rect 463 -121 497 -105
rect 463 -313 497 -297
rect -465 -381 -449 -347
rect -415 -381 -399 -347
rect -273 -381 -257 -347
rect -223 -381 -207 -347
rect -81 -381 -65 -347
rect -31 -381 -15 -347
rect 111 -381 127 -347
rect 161 -381 177 -347
rect 303 -381 319 -347
rect 353 -381 369 -347
rect -465 -489 -449 -455
rect -415 -489 -399 -455
rect -273 -489 -257 -455
rect -223 -489 -207 -455
rect -81 -489 -65 -455
rect -31 -489 -15 -455
rect 111 -489 127 -455
rect 161 -489 177 -455
rect 303 -489 319 -455
rect 353 -489 369 -455
rect -497 -539 -463 -523
rect -497 -731 -463 -715
rect -401 -539 -367 -523
rect -401 -731 -367 -715
rect -305 -539 -271 -523
rect -305 -731 -271 -715
rect -209 -539 -175 -523
rect -209 -731 -175 -715
rect -113 -539 -79 -523
rect -113 -731 -79 -715
rect -17 -539 17 -523
rect -17 -731 17 -715
rect 79 -539 113 -523
rect 79 -731 113 -715
rect 175 -539 209 -523
rect 175 -731 209 -715
rect 271 -539 305 -523
rect 271 -731 305 -715
rect 367 -539 401 -523
rect 367 -731 401 -715
rect 463 -539 497 -523
rect 463 -731 497 -715
rect -369 -799 -353 -765
rect -319 -799 -303 -765
rect -177 -799 -161 -765
rect -127 -799 -111 -765
rect 15 -799 31 -765
rect 65 -799 81 -765
rect 207 -799 223 -765
rect 257 -799 273 -765
rect 399 -799 415 -765
rect 449 -799 465 -765
rect -369 -907 -353 -873
rect -319 -907 -303 -873
rect -177 -907 -161 -873
rect -127 -907 -111 -873
rect 15 -907 31 -873
rect 65 -907 81 -873
rect 207 -907 223 -873
rect 257 -907 273 -873
rect 399 -907 415 -873
rect 449 -907 465 -873
rect -497 -957 -463 -941
rect -497 -1149 -463 -1133
rect -401 -957 -367 -941
rect -401 -1149 -367 -1133
rect -305 -957 -271 -941
rect -305 -1149 -271 -1133
rect -209 -957 -175 -941
rect -209 -1149 -175 -1133
rect -113 -957 -79 -941
rect -113 -1149 -79 -1133
rect -17 -957 17 -941
rect -17 -1149 17 -1133
rect 79 -957 113 -941
rect 79 -1149 113 -1133
rect 175 -957 209 -941
rect 175 -1149 209 -1133
rect 271 -957 305 -941
rect 271 -1149 305 -1133
rect 367 -957 401 -941
rect 367 -1149 401 -1133
rect 463 -957 497 -941
rect 463 -1149 497 -1133
rect -465 -1217 -449 -1183
rect -415 -1217 -399 -1183
rect -273 -1217 -257 -1183
rect -223 -1217 -207 -1183
rect -81 -1217 -65 -1183
rect -31 -1217 -15 -1183
rect 111 -1217 127 -1183
rect 161 -1217 177 -1183
rect 303 -1217 319 -1183
rect 353 -1217 369 -1183
rect -611 -1285 -577 -1223
rect 577 -1285 611 -1223
rect -611 -1319 -515 -1285
rect 515 -1319 611 -1285
<< viali >>
rect -449 1183 -415 1217
rect -257 1183 -223 1217
rect -65 1183 -31 1217
rect 127 1183 161 1217
rect 319 1183 353 1217
rect -497 957 -463 1133
rect -401 957 -367 1133
rect -305 957 -271 1133
rect -209 957 -175 1133
rect -113 957 -79 1133
rect -17 957 17 1133
rect 79 957 113 1133
rect 175 957 209 1133
rect 271 957 305 1133
rect 367 957 401 1133
rect 463 957 497 1133
rect -353 873 -319 907
rect -161 873 -127 907
rect 31 873 65 907
rect 223 873 257 907
rect 415 873 449 907
rect -353 765 -319 799
rect -161 765 -127 799
rect 31 765 65 799
rect 223 765 257 799
rect 415 765 449 799
rect -497 539 -463 715
rect -401 539 -367 715
rect -305 539 -271 715
rect -209 539 -175 715
rect -113 539 -79 715
rect -17 539 17 715
rect 79 539 113 715
rect 175 539 209 715
rect 271 539 305 715
rect 367 539 401 715
rect 463 539 497 715
rect -449 455 -415 489
rect -257 455 -223 489
rect -65 455 -31 489
rect 127 455 161 489
rect 319 455 353 489
rect -449 347 -415 381
rect -257 347 -223 381
rect -65 347 -31 381
rect 127 347 161 381
rect 319 347 353 381
rect -497 121 -463 297
rect -401 121 -367 297
rect -305 121 -271 297
rect -209 121 -175 297
rect -113 121 -79 297
rect -17 121 17 297
rect 79 121 113 297
rect 175 121 209 297
rect 271 121 305 297
rect 367 121 401 297
rect 463 121 497 297
rect -353 37 -319 71
rect -161 37 -127 71
rect 31 37 65 71
rect 223 37 257 71
rect 415 37 449 71
rect -353 -71 -319 -37
rect -161 -71 -127 -37
rect 31 -71 65 -37
rect 223 -71 257 -37
rect 415 -71 449 -37
rect -497 -297 -463 -121
rect -401 -297 -367 -121
rect -305 -297 -271 -121
rect -209 -297 -175 -121
rect -113 -297 -79 -121
rect -17 -297 17 -121
rect 79 -297 113 -121
rect 175 -297 209 -121
rect 271 -297 305 -121
rect 367 -297 401 -121
rect 463 -297 497 -121
rect -449 -381 -415 -347
rect -257 -381 -223 -347
rect -65 -381 -31 -347
rect 127 -381 161 -347
rect 319 -381 353 -347
rect -449 -489 -415 -455
rect -257 -489 -223 -455
rect -65 -489 -31 -455
rect 127 -489 161 -455
rect 319 -489 353 -455
rect -497 -715 -463 -539
rect -401 -715 -367 -539
rect -305 -715 -271 -539
rect -209 -715 -175 -539
rect -113 -715 -79 -539
rect -17 -715 17 -539
rect 79 -715 113 -539
rect 175 -715 209 -539
rect 271 -715 305 -539
rect 367 -715 401 -539
rect 463 -715 497 -539
rect -353 -799 -319 -765
rect -161 -799 -127 -765
rect 31 -799 65 -765
rect 223 -799 257 -765
rect 415 -799 449 -765
rect -353 -907 -319 -873
rect -161 -907 -127 -873
rect 31 -907 65 -873
rect 223 -907 257 -873
rect 415 -907 449 -873
rect -497 -1133 -463 -957
rect -401 -1133 -367 -957
rect -305 -1133 -271 -957
rect -209 -1133 -175 -957
rect -113 -1133 -79 -957
rect -17 -1133 17 -957
rect 79 -1133 113 -957
rect 175 -1133 209 -957
rect 271 -1133 305 -957
rect 367 -1133 401 -957
rect 463 -1133 497 -957
rect -449 -1217 -415 -1183
rect -257 -1217 -223 -1183
rect -65 -1217 -31 -1183
rect 127 -1217 161 -1183
rect 319 -1217 353 -1183
<< metal1 >>
rect -461 1217 -403 1223
rect -461 1183 -449 1217
rect -415 1183 -403 1217
rect -461 1177 -403 1183
rect -269 1217 -211 1223
rect -269 1183 -257 1217
rect -223 1183 -211 1217
rect -269 1177 -211 1183
rect -77 1217 -19 1223
rect -77 1183 -65 1217
rect -31 1183 -19 1217
rect -77 1177 -19 1183
rect 115 1217 173 1223
rect 115 1183 127 1217
rect 161 1183 173 1217
rect 115 1177 173 1183
rect 307 1217 365 1223
rect 307 1183 319 1217
rect 353 1183 365 1217
rect 307 1177 365 1183
rect -503 1133 -457 1145
rect -503 957 -497 1133
rect -463 957 -457 1133
rect -503 945 -457 957
rect -407 1133 -361 1145
rect -407 957 -401 1133
rect -367 957 -361 1133
rect -407 945 -361 957
rect -311 1133 -265 1145
rect -311 957 -305 1133
rect -271 957 -265 1133
rect -311 945 -265 957
rect -215 1133 -169 1145
rect -215 957 -209 1133
rect -175 957 -169 1133
rect -215 945 -169 957
rect -119 1133 -73 1145
rect -119 957 -113 1133
rect -79 957 -73 1133
rect -119 945 -73 957
rect -23 1133 23 1145
rect -23 957 -17 1133
rect 17 957 23 1133
rect -23 945 23 957
rect 73 1133 119 1145
rect 73 957 79 1133
rect 113 957 119 1133
rect 73 945 119 957
rect 169 1133 215 1145
rect 169 957 175 1133
rect 209 957 215 1133
rect 169 945 215 957
rect 265 1133 311 1145
rect 265 957 271 1133
rect 305 957 311 1133
rect 265 945 311 957
rect 361 1133 407 1145
rect 361 957 367 1133
rect 401 957 407 1133
rect 361 945 407 957
rect 457 1133 503 1145
rect 457 957 463 1133
rect 497 957 503 1133
rect 457 945 503 957
rect -365 907 -307 913
rect -365 873 -353 907
rect -319 873 -307 907
rect -365 867 -307 873
rect -173 907 -115 913
rect -173 873 -161 907
rect -127 873 -115 907
rect -173 867 -115 873
rect 19 907 77 913
rect 19 873 31 907
rect 65 873 77 907
rect 19 867 77 873
rect 211 907 269 913
rect 211 873 223 907
rect 257 873 269 907
rect 211 867 269 873
rect 403 907 461 913
rect 403 873 415 907
rect 449 873 461 907
rect 403 867 461 873
rect -365 799 -307 805
rect -365 765 -353 799
rect -319 765 -307 799
rect -365 759 -307 765
rect -173 799 -115 805
rect -173 765 -161 799
rect -127 765 -115 799
rect -173 759 -115 765
rect 19 799 77 805
rect 19 765 31 799
rect 65 765 77 799
rect 19 759 77 765
rect 211 799 269 805
rect 211 765 223 799
rect 257 765 269 799
rect 211 759 269 765
rect 403 799 461 805
rect 403 765 415 799
rect 449 765 461 799
rect 403 759 461 765
rect -503 715 -457 727
rect -503 539 -497 715
rect -463 539 -457 715
rect -503 527 -457 539
rect -407 715 -361 727
rect -407 539 -401 715
rect -367 539 -361 715
rect -407 527 -361 539
rect -311 715 -265 727
rect -311 539 -305 715
rect -271 539 -265 715
rect -311 527 -265 539
rect -215 715 -169 727
rect -215 539 -209 715
rect -175 539 -169 715
rect -215 527 -169 539
rect -119 715 -73 727
rect -119 539 -113 715
rect -79 539 -73 715
rect -119 527 -73 539
rect -23 715 23 727
rect -23 539 -17 715
rect 17 539 23 715
rect -23 527 23 539
rect 73 715 119 727
rect 73 539 79 715
rect 113 539 119 715
rect 73 527 119 539
rect 169 715 215 727
rect 169 539 175 715
rect 209 539 215 715
rect 169 527 215 539
rect 265 715 311 727
rect 265 539 271 715
rect 305 539 311 715
rect 265 527 311 539
rect 361 715 407 727
rect 361 539 367 715
rect 401 539 407 715
rect 361 527 407 539
rect 457 715 503 727
rect 457 539 463 715
rect 497 539 503 715
rect 457 527 503 539
rect -461 489 -403 495
rect -461 455 -449 489
rect -415 455 -403 489
rect -461 449 -403 455
rect -269 489 -211 495
rect -269 455 -257 489
rect -223 455 -211 489
rect -269 449 -211 455
rect -77 489 -19 495
rect -77 455 -65 489
rect -31 455 -19 489
rect -77 449 -19 455
rect 115 489 173 495
rect 115 455 127 489
rect 161 455 173 489
rect 115 449 173 455
rect 307 489 365 495
rect 307 455 319 489
rect 353 455 365 489
rect 307 449 365 455
rect -461 381 -403 387
rect -461 347 -449 381
rect -415 347 -403 381
rect -461 341 -403 347
rect -269 381 -211 387
rect -269 347 -257 381
rect -223 347 -211 381
rect -269 341 -211 347
rect -77 381 -19 387
rect -77 347 -65 381
rect -31 347 -19 381
rect -77 341 -19 347
rect 115 381 173 387
rect 115 347 127 381
rect 161 347 173 381
rect 115 341 173 347
rect 307 381 365 387
rect 307 347 319 381
rect 353 347 365 381
rect 307 341 365 347
rect -503 297 -457 309
rect -503 121 -497 297
rect -463 121 -457 297
rect -503 109 -457 121
rect -407 297 -361 309
rect -407 121 -401 297
rect -367 121 -361 297
rect -407 109 -361 121
rect -311 297 -265 309
rect -311 121 -305 297
rect -271 121 -265 297
rect -311 109 -265 121
rect -215 297 -169 309
rect -215 121 -209 297
rect -175 121 -169 297
rect -215 109 -169 121
rect -119 297 -73 309
rect -119 121 -113 297
rect -79 121 -73 297
rect -119 109 -73 121
rect -23 297 23 309
rect -23 121 -17 297
rect 17 121 23 297
rect -23 109 23 121
rect 73 297 119 309
rect 73 121 79 297
rect 113 121 119 297
rect 73 109 119 121
rect 169 297 215 309
rect 169 121 175 297
rect 209 121 215 297
rect 169 109 215 121
rect 265 297 311 309
rect 265 121 271 297
rect 305 121 311 297
rect 265 109 311 121
rect 361 297 407 309
rect 361 121 367 297
rect 401 121 407 297
rect 361 109 407 121
rect 457 297 503 309
rect 457 121 463 297
rect 497 121 503 297
rect 457 109 503 121
rect -365 71 -307 77
rect -365 37 -353 71
rect -319 37 -307 71
rect -365 31 -307 37
rect -173 71 -115 77
rect -173 37 -161 71
rect -127 37 -115 71
rect -173 31 -115 37
rect 19 71 77 77
rect 19 37 31 71
rect 65 37 77 71
rect 19 31 77 37
rect 211 71 269 77
rect 211 37 223 71
rect 257 37 269 71
rect 211 31 269 37
rect 403 71 461 77
rect 403 37 415 71
rect 449 37 461 71
rect 403 31 461 37
rect -365 -37 -307 -31
rect -365 -71 -353 -37
rect -319 -71 -307 -37
rect -365 -77 -307 -71
rect -173 -37 -115 -31
rect -173 -71 -161 -37
rect -127 -71 -115 -37
rect -173 -77 -115 -71
rect 19 -37 77 -31
rect 19 -71 31 -37
rect 65 -71 77 -37
rect 19 -77 77 -71
rect 211 -37 269 -31
rect 211 -71 223 -37
rect 257 -71 269 -37
rect 211 -77 269 -71
rect 403 -37 461 -31
rect 403 -71 415 -37
rect 449 -71 461 -37
rect 403 -77 461 -71
rect -503 -121 -457 -109
rect -503 -297 -497 -121
rect -463 -297 -457 -121
rect -503 -309 -457 -297
rect -407 -121 -361 -109
rect -407 -297 -401 -121
rect -367 -297 -361 -121
rect -407 -309 -361 -297
rect -311 -121 -265 -109
rect -311 -297 -305 -121
rect -271 -297 -265 -121
rect -311 -309 -265 -297
rect -215 -121 -169 -109
rect -215 -297 -209 -121
rect -175 -297 -169 -121
rect -215 -309 -169 -297
rect -119 -121 -73 -109
rect -119 -297 -113 -121
rect -79 -297 -73 -121
rect -119 -309 -73 -297
rect -23 -121 23 -109
rect -23 -297 -17 -121
rect 17 -297 23 -121
rect -23 -309 23 -297
rect 73 -121 119 -109
rect 73 -297 79 -121
rect 113 -297 119 -121
rect 73 -309 119 -297
rect 169 -121 215 -109
rect 169 -297 175 -121
rect 209 -297 215 -121
rect 169 -309 215 -297
rect 265 -121 311 -109
rect 265 -297 271 -121
rect 305 -297 311 -121
rect 265 -309 311 -297
rect 361 -121 407 -109
rect 361 -297 367 -121
rect 401 -297 407 -121
rect 361 -309 407 -297
rect 457 -121 503 -109
rect 457 -297 463 -121
rect 497 -297 503 -121
rect 457 -309 503 -297
rect -461 -347 -403 -341
rect -461 -381 -449 -347
rect -415 -381 -403 -347
rect -461 -387 -403 -381
rect -269 -347 -211 -341
rect -269 -381 -257 -347
rect -223 -381 -211 -347
rect -269 -387 -211 -381
rect -77 -347 -19 -341
rect -77 -381 -65 -347
rect -31 -381 -19 -347
rect -77 -387 -19 -381
rect 115 -347 173 -341
rect 115 -381 127 -347
rect 161 -381 173 -347
rect 115 -387 173 -381
rect 307 -347 365 -341
rect 307 -381 319 -347
rect 353 -381 365 -347
rect 307 -387 365 -381
rect -461 -455 -403 -449
rect -461 -489 -449 -455
rect -415 -489 -403 -455
rect -461 -495 -403 -489
rect -269 -455 -211 -449
rect -269 -489 -257 -455
rect -223 -489 -211 -455
rect -269 -495 -211 -489
rect -77 -455 -19 -449
rect -77 -489 -65 -455
rect -31 -489 -19 -455
rect -77 -495 -19 -489
rect 115 -455 173 -449
rect 115 -489 127 -455
rect 161 -489 173 -455
rect 115 -495 173 -489
rect 307 -455 365 -449
rect 307 -489 319 -455
rect 353 -489 365 -455
rect 307 -495 365 -489
rect -503 -539 -457 -527
rect -503 -715 -497 -539
rect -463 -715 -457 -539
rect -503 -727 -457 -715
rect -407 -539 -361 -527
rect -407 -715 -401 -539
rect -367 -715 -361 -539
rect -407 -727 -361 -715
rect -311 -539 -265 -527
rect -311 -715 -305 -539
rect -271 -715 -265 -539
rect -311 -727 -265 -715
rect -215 -539 -169 -527
rect -215 -715 -209 -539
rect -175 -715 -169 -539
rect -215 -727 -169 -715
rect -119 -539 -73 -527
rect -119 -715 -113 -539
rect -79 -715 -73 -539
rect -119 -727 -73 -715
rect -23 -539 23 -527
rect -23 -715 -17 -539
rect 17 -715 23 -539
rect -23 -727 23 -715
rect 73 -539 119 -527
rect 73 -715 79 -539
rect 113 -715 119 -539
rect 73 -727 119 -715
rect 169 -539 215 -527
rect 169 -715 175 -539
rect 209 -715 215 -539
rect 169 -727 215 -715
rect 265 -539 311 -527
rect 265 -715 271 -539
rect 305 -715 311 -539
rect 265 -727 311 -715
rect 361 -539 407 -527
rect 361 -715 367 -539
rect 401 -715 407 -539
rect 361 -727 407 -715
rect 457 -539 503 -527
rect 457 -715 463 -539
rect 497 -715 503 -539
rect 457 -727 503 -715
rect -365 -765 -307 -759
rect -365 -799 -353 -765
rect -319 -799 -307 -765
rect -365 -805 -307 -799
rect -173 -765 -115 -759
rect -173 -799 -161 -765
rect -127 -799 -115 -765
rect -173 -805 -115 -799
rect 19 -765 77 -759
rect 19 -799 31 -765
rect 65 -799 77 -765
rect 19 -805 77 -799
rect 211 -765 269 -759
rect 211 -799 223 -765
rect 257 -799 269 -765
rect 211 -805 269 -799
rect 403 -765 461 -759
rect 403 -799 415 -765
rect 449 -799 461 -765
rect 403 -805 461 -799
rect -365 -873 -307 -867
rect -365 -907 -353 -873
rect -319 -907 -307 -873
rect -365 -913 -307 -907
rect -173 -873 -115 -867
rect -173 -907 -161 -873
rect -127 -907 -115 -873
rect -173 -913 -115 -907
rect 19 -873 77 -867
rect 19 -907 31 -873
rect 65 -907 77 -873
rect 19 -913 77 -907
rect 211 -873 269 -867
rect 211 -907 223 -873
rect 257 -907 269 -873
rect 211 -913 269 -907
rect 403 -873 461 -867
rect 403 -907 415 -873
rect 449 -907 461 -873
rect 403 -913 461 -907
rect -503 -957 -457 -945
rect -503 -1133 -497 -957
rect -463 -1133 -457 -957
rect -503 -1145 -457 -1133
rect -407 -957 -361 -945
rect -407 -1133 -401 -957
rect -367 -1133 -361 -957
rect -407 -1145 -361 -1133
rect -311 -957 -265 -945
rect -311 -1133 -305 -957
rect -271 -1133 -265 -957
rect -311 -1145 -265 -1133
rect -215 -957 -169 -945
rect -215 -1133 -209 -957
rect -175 -1133 -169 -957
rect -215 -1145 -169 -1133
rect -119 -957 -73 -945
rect -119 -1133 -113 -957
rect -79 -1133 -73 -957
rect -119 -1145 -73 -1133
rect -23 -957 23 -945
rect -23 -1133 -17 -957
rect 17 -1133 23 -957
rect -23 -1145 23 -1133
rect 73 -957 119 -945
rect 73 -1133 79 -957
rect 113 -1133 119 -957
rect 73 -1145 119 -1133
rect 169 -957 215 -945
rect 169 -1133 175 -957
rect 209 -1133 215 -957
rect 169 -1145 215 -1133
rect 265 -957 311 -945
rect 265 -1133 271 -957
rect 305 -1133 311 -957
rect 265 -1145 311 -1133
rect 361 -957 407 -945
rect 361 -1133 367 -957
rect 401 -1133 407 -957
rect 361 -1145 407 -1133
rect 457 -957 503 -945
rect 457 -1133 463 -957
rect 497 -1133 503 -957
rect 457 -1145 503 -1133
rect -461 -1183 -403 -1177
rect -461 -1217 -449 -1183
rect -415 -1217 -403 -1183
rect -461 -1223 -403 -1217
rect -269 -1183 -211 -1177
rect -269 -1217 -257 -1183
rect -223 -1217 -211 -1183
rect -269 -1223 -211 -1217
rect -77 -1183 -19 -1177
rect -77 -1217 -65 -1183
rect -31 -1217 -19 -1183
rect -77 -1223 -19 -1217
rect 115 -1183 173 -1177
rect 115 -1217 127 -1183
rect 161 -1217 173 -1183
rect 115 -1223 173 -1217
rect 307 -1183 365 -1177
rect 307 -1217 319 -1183
rect 353 -1217 365 -1183
rect 307 -1223 365 -1217
<< properties >>
string FIXED_BBOX -594 -1302 594 1302
string gencell sky130_fd_pr__nfet_01v8_lvt
string library sky130
string parameters w 1.0 l 0.15 m 6 nf 10 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
