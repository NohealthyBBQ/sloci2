magic
tech sky130A
magscale 1 2
timestamp 1662976792
<< pwell >>
rect 53403 -7310 53408 -7308
<< ndiff >>
rect 53403 -7310 53408 -7308
<< locali >>
rect 48302 -6542 48426 -6396
rect 51418 -6516 51882 -6426
rect 64120 -6540 64294 -6402
rect 68132 -6542 68246 -6400
<< viali >>
rect 48286 -5236 48458 -5178
rect 49920 -5280 66568 -5188
rect 68070 -5236 68242 -5178
rect 48274 -7764 48446 -7706
rect 49940 -7756 66588 -7664
rect 68120 -7768 68292 -7710
<< metal1 >>
rect 48274 -5178 48470 -5172
rect 47250 -6264 47260 -5190
rect 47620 -6264 47630 -5190
rect 48274 -5236 48286 -5178
rect 48458 -5236 48470 -5178
rect 68058 -5178 68254 -5172
rect 48274 -5242 48470 -5236
rect 49908 -5188 66580 -5182
rect 49908 -5280 49920 -5188
rect 66568 -5280 66580 -5188
rect 68058 -5236 68070 -5178
rect 68242 -5236 68254 -5178
rect 68058 -5242 68254 -5236
rect 49908 -5286 66580 -5280
rect 48190 -5686 48550 -5300
rect 48188 -6296 48550 -5686
rect 49880 -5400 66630 -5370
rect 49880 -5680 49910 -5400
rect 50077 -5494 50087 -5442
rect 50139 -5494 50149 -5442
rect 50267 -5493 50277 -5441
rect 50329 -5493 50339 -5441
rect 50460 -5496 50470 -5444
rect 50522 -5496 50532 -5444
rect 50652 -5491 50662 -5439
rect 50714 -5491 50724 -5439
rect 50844 -5495 50854 -5443
rect 50906 -5495 50916 -5443
rect 51036 -5490 51046 -5438
rect 51098 -5490 51108 -5438
rect 51228 -5491 51238 -5439
rect 51290 -5491 51300 -5439
rect 51418 -5490 51428 -5438
rect 51480 -5490 51490 -5438
rect 51612 -5501 51622 -5449
rect 51674 -5501 51684 -5449
rect 51801 -5499 51811 -5447
rect 51863 -5499 51873 -5447
rect 51991 -5499 52001 -5447
rect 52053 -5499 52063 -5447
rect 52190 -5500 52200 -5448
rect 52252 -5500 52262 -5448
rect 52382 -5499 52392 -5447
rect 52444 -5499 52454 -5447
rect 52572 -5500 52582 -5448
rect 52634 -5500 52644 -5448
rect 52764 -5493 52774 -5441
rect 52826 -5493 52836 -5441
rect 52956 -5495 52966 -5443
rect 53018 -5495 53028 -5443
rect 53149 -5494 53159 -5442
rect 53211 -5494 53221 -5442
rect 53341 -5492 53351 -5440
rect 53403 -5492 53413 -5440
rect 53532 -5492 53542 -5440
rect 53594 -5492 53604 -5440
rect 53726 -5497 53736 -5445
rect 53788 -5497 53798 -5445
rect 53917 -5493 53927 -5441
rect 53979 -5493 53989 -5441
rect 54109 -5489 54119 -5437
rect 54171 -5489 54181 -5437
rect 54302 -5493 54312 -5441
rect 54364 -5493 54374 -5441
rect 54494 -5493 54504 -5441
rect 54556 -5493 54566 -5441
rect 54687 -5494 54697 -5442
rect 54749 -5494 54759 -5442
rect 54879 -5492 54889 -5440
rect 54941 -5492 54951 -5440
rect 55070 -5491 55080 -5439
rect 55132 -5491 55142 -5439
rect 55261 -5490 55271 -5438
rect 55323 -5490 55333 -5438
rect 55454 -5490 55464 -5438
rect 55516 -5490 55526 -5438
rect 55645 -5499 55655 -5447
rect 55707 -5499 55717 -5447
rect 55836 -5500 55846 -5448
rect 55898 -5500 55908 -5448
rect 56026 -5501 56036 -5449
rect 56088 -5501 56098 -5449
rect 56220 -5505 56230 -5453
rect 56282 -5505 56292 -5453
rect 56412 -5507 56422 -5455
rect 56474 -5507 56484 -5455
rect 56606 -5506 56616 -5454
rect 56668 -5506 56678 -5454
rect 56798 -5503 56808 -5451
rect 56860 -5503 56870 -5451
rect 56987 -5500 56997 -5448
rect 57049 -5500 57059 -5448
rect 57181 -5498 57191 -5446
rect 57243 -5498 57253 -5446
rect 57374 -5499 57384 -5447
rect 57436 -5499 57446 -5447
rect 57567 -5500 57577 -5448
rect 57629 -5500 57639 -5448
rect 57756 -5500 57766 -5448
rect 57818 -5500 57828 -5448
rect 57949 -5500 57959 -5448
rect 58011 -5500 58021 -5448
rect 58141 -5500 58151 -5448
rect 58203 -5500 58213 -5448
rect 58332 -5500 58342 -5448
rect 58394 -5500 58404 -5448
rect 58525 -5500 58535 -5448
rect 58587 -5500 58597 -5448
rect 58716 -5499 58726 -5447
rect 58778 -5499 58788 -5447
rect 58911 -5500 58921 -5448
rect 58973 -5500 58983 -5448
rect 59100 -5500 59110 -5448
rect 59162 -5500 59172 -5448
rect 59293 -5500 59303 -5448
rect 59355 -5500 59365 -5448
rect 59485 -5500 59495 -5448
rect 59547 -5500 59557 -5448
rect 59676 -5500 59686 -5448
rect 59738 -5500 59748 -5448
rect 59868 -5500 59878 -5448
rect 59930 -5500 59940 -5448
rect 60061 -5500 60071 -5448
rect 60123 -5500 60133 -5448
rect 60250 -5501 60260 -5449
rect 60312 -5501 60322 -5449
rect 60444 -5500 60454 -5448
rect 60506 -5500 60516 -5448
rect 60635 -5500 60645 -5448
rect 60697 -5500 60707 -5448
rect 60828 -5500 60838 -5448
rect 60890 -5500 60900 -5448
rect 61020 -5500 61030 -5448
rect 61082 -5500 61092 -5448
rect 61212 -5501 61222 -5449
rect 61274 -5501 61284 -5449
rect 61405 -5499 61415 -5447
rect 61467 -5499 61477 -5447
rect 61595 -5499 61605 -5447
rect 61657 -5499 61667 -5447
rect 61788 -5501 61798 -5449
rect 61850 -5501 61860 -5449
rect 61980 -5500 61990 -5448
rect 62042 -5500 62052 -5448
rect 62173 -5499 62183 -5447
rect 62235 -5499 62245 -5447
rect 62364 -5499 62374 -5447
rect 62426 -5499 62436 -5447
rect 62556 -5500 62566 -5448
rect 62618 -5500 62628 -5448
rect 62747 -5500 62757 -5448
rect 62809 -5500 62819 -5448
rect 62939 -5500 62949 -5448
rect 63001 -5500 63011 -5448
rect 63133 -5499 63143 -5447
rect 63195 -5499 63205 -5447
rect 63325 -5500 63335 -5448
rect 63387 -5500 63397 -5448
rect 63515 -5501 63525 -5449
rect 63577 -5501 63587 -5449
rect 63706 -5502 63716 -5450
rect 63768 -5502 63778 -5450
rect 63899 -5500 63909 -5448
rect 63961 -5500 63971 -5448
rect 64092 -5499 64102 -5447
rect 64154 -5499 64164 -5447
rect 64285 -5500 64295 -5448
rect 64347 -5500 64357 -5448
rect 64476 -5500 64486 -5448
rect 64538 -5500 64548 -5448
rect 64667 -5500 64677 -5448
rect 64729 -5500 64739 -5448
rect 64860 -5500 64870 -5448
rect 64922 -5500 64932 -5448
rect 65053 -5500 65063 -5448
rect 65115 -5500 65125 -5448
rect 65244 -5500 65254 -5448
rect 65306 -5500 65316 -5448
rect 65435 -5499 65445 -5447
rect 65497 -5499 65507 -5447
rect 65626 -5499 65636 -5447
rect 65688 -5499 65698 -5447
rect 65819 -5500 65829 -5448
rect 65881 -5500 65891 -5448
rect 66013 -5500 66023 -5448
rect 66075 -5500 66085 -5448
rect 66201 -5501 66211 -5449
rect 66263 -5501 66273 -5449
rect 66395 -5509 66405 -5457
rect 66457 -5509 66467 -5457
rect 49981 -5637 49991 -5585
rect 50043 -5637 50053 -5585
rect 50172 -5639 50182 -5587
rect 50234 -5639 50244 -5587
rect 50364 -5638 50374 -5586
rect 50426 -5638 50436 -5586
rect 50556 -5641 50566 -5589
rect 50618 -5641 50628 -5589
rect 50750 -5640 50760 -5588
rect 50812 -5640 50822 -5588
rect 50940 -5640 50950 -5588
rect 51002 -5640 51012 -5588
rect 51135 -5638 51145 -5586
rect 51197 -5638 51207 -5586
rect 51326 -5637 51336 -5585
rect 51388 -5637 51398 -5585
rect 51521 -5639 51531 -5587
rect 51583 -5639 51593 -5587
rect 51711 -5639 51721 -5587
rect 51773 -5639 51783 -5587
rect 51901 -5638 51911 -5586
rect 51963 -5638 51973 -5586
rect 52094 -5637 52104 -5585
rect 52156 -5637 52166 -5585
rect 52285 -5637 52295 -5585
rect 52347 -5637 52357 -5585
rect 52481 -5639 52491 -5587
rect 52543 -5639 52553 -5587
rect 52670 -5639 52680 -5587
rect 52732 -5639 52742 -5587
rect 52864 -5639 52874 -5587
rect 52926 -5639 52936 -5587
rect 53053 -5639 53063 -5587
rect 53115 -5639 53125 -5587
rect 53245 -5640 53255 -5588
rect 53307 -5640 53317 -5588
rect 53438 -5640 53448 -5588
rect 53500 -5640 53510 -5588
rect 53629 -5640 53639 -5588
rect 53691 -5640 53701 -5588
rect 53821 -5639 53831 -5587
rect 53883 -5639 53893 -5587
rect 54013 -5640 54023 -5588
rect 54075 -5640 54085 -5588
rect 54206 -5640 54216 -5588
rect 54268 -5640 54278 -5588
rect 54397 -5640 54407 -5588
rect 54459 -5640 54469 -5588
rect 54589 -5639 54599 -5587
rect 54651 -5639 54661 -5587
rect 54782 -5640 54792 -5588
rect 54844 -5640 54854 -5588
rect 54974 -5640 54984 -5588
rect 55036 -5640 55046 -5588
rect 55165 -5640 55175 -5588
rect 55227 -5640 55237 -5588
rect 55356 -5640 55366 -5588
rect 55418 -5640 55428 -5588
rect 55548 -5640 55558 -5588
rect 55610 -5640 55620 -5588
rect 55741 -5639 55751 -5587
rect 55803 -5639 55813 -5587
rect 55932 -5639 55942 -5587
rect 55994 -5639 56004 -5587
rect 56126 -5640 56136 -5588
rect 56188 -5640 56198 -5588
rect 56318 -5640 56328 -5588
rect 56380 -5640 56390 -5588
rect 56510 -5640 56520 -5588
rect 56572 -5640 56582 -5588
rect 56702 -5640 56712 -5588
rect 56764 -5640 56774 -5588
rect 56894 -5640 56904 -5588
rect 56956 -5640 56966 -5588
rect 57086 -5640 57096 -5588
rect 57148 -5640 57158 -5588
rect 57278 -5640 57288 -5588
rect 57340 -5640 57350 -5588
rect 57469 -5640 57479 -5588
rect 57531 -5640 57541 -5588
rect 57661 -5640 57671 -5588
rect 57723 -5640 57733 -5588
rect 57854 -5640 57864 -5588
rect 57916 -5640 57926 -5588
rect 58046 -5640 58056 -5588
rect 58108 -5640 58118 -5588
rect 58238 -5640 58248 -5588
rect 58300 -5640 58310 -5588
rect 58429 -5640 58439 -5588
rect 58491 -5640 58501 -5588
rect 58621 -5640 58631 -5588
rect 58683 -5640 58693 -5588
rect 58812 -5640 58822 -5588
rect 58874 -5640 58884 -5588
rect 59003 -5640 59013 -5588
rect 59065 -5640 59075 -5588
rect 59197 -5640 59207 -5588
rect 59259 -5640 59269 -5588
rect 59389 -5640 59399 -5588
rect 59451 -5640 59461 -5588
rect 59582 -5639 59592 -5587
rect 59644 -5639 59654 -5587
rect 59773 -5640 59783 -5588
rect 59835 -5640 59845 -5588
rect 59965 -5640 59975 -5588
rect 60027 -5640 60037 -5588
rect 60158 -5640 60168 -5588
rect 60220 -5640 60230 -5588
rect 60350 -5640 60360 -5588
rect 60412 -5640 60422 -5588
rect 60543 -5639 60553 -5587
rect 60605 -5639 60615 -5587
rect 60734 -5640 60744 -5588
rect 60796 -5640 60806 -5588
rect 60926 -5640 60936 -5588
rect 60988 -5640 60998 -5588
rect 61117 -5640 61127 -5588
rect 61179 -5640 61189 -5588
rect 61309 -5640 61319 -5588
rect 61371 -5640 61381 -5588
rect 61501 -5640 61511 -5588
rect 61563 -5640 61573 -5588
rect 61694 -5640 61704 -5588
rect 61756 -5640 61766 -5588
rect 61885 -5640 61895 -5588
rect 61947 -5640 61957 -5588
rect 62077 -5640 62087 -5588
rect 62139 -5640 62149 -5588
rect 62269 -5639 62279 -5587
rect 62331 -5639 62341 -5587
rect 62461 -5640 62471 -5588
rect 62523 -5640 62533 -5588
rect 62651 -5640 62661 -5588
rect 62713 -5640 62723 -5588
rect 62845 -5640 62855 -5588
rect 62907 -5640 62917 -5588
rect 63037 -5639 63047 -5587
rect 63099 -5639 63109 -5587
rect 63228 -5640 63238 -5588
rect 63290 -5640 63300 -5588
rect 63421 -5640 63431 -5588
rect 63483 -5640 63493 -5588
rect 63612 -5639 63622 -5587
rect 63674 -5639 63684 -5587
rect 63804 -5640 63814 -5588
rect 63866 -5640 63876 -5588
rect 63995 -5640 64005 -5588
rect 64057 -5640 64067 -5588
rect 64189 -5639 64199 -5587
rect 64251 -5639 64261 -5587
rect 64380 -5640 64390 -5588
rect 64442 -5640 64452 -5588
rect 64572 -5640 64582 -5588
rect 64634 -5640 64644 -5588
rect 64764 -5640 64774 -5588
rect 64826 -5640 64836 -5588
rect 64956 -5640 64966 -5588
rect 65018 -5640 65028 -5588
rect 65149 -5640 65159 -5588
rect 65211 -5640 65221 -5588
rect 65340 -5640 65350 -5588
rect 65402 -5640 65412 -5588
rect 65533 -5639 65543 -5587
rect 65595 -5639 65605 -5587
rect 65724 -5640 65734 -5588
rect 65786 -5640 65796 -5588
rect 65917 -5640 65927 -5588
rect 65979 -5640 65989 -5588
rect 66108 -5640 66118 -5588
rect 66170 -5640 66180 -5588
rect 66299 -5638 66309 -5586
rect 66361 -5638 66371 -5586
rect 66494 -5640 66504 -5588
rect 66556 -5640 66566 -5588
rect 66600 -5680 66630 -5400
rect 49880 -5710 66630 -5680
rect 68000 -5710 68374 -5302
rect 51860 -6020 57940 -5990
rect 49420 -6126 49430 -6074
rect 49482 -6126 49492 -6074
rect 51860 -6300 51890 -6020
rect 52037 -6123 52047 -6071
rect 52099 -6123 52109 -6071
rect 52227 -6122 52237 -6070
rect 52289 -6122 52299 -6070
rect 52419 -6121 52429 -6069
rect 52481 -6121 52491 -6069
rect 52610 -6121 52620 -6069
rect 52672 -6121 52682 -6069
rect 52804 -6121 52814 -6069
rect 52866 -6121 52876 -6069
rect 52994 -6122 53004 -6070
rect 53056 -6122 53066 -6070
rect 53188 -6121 53198 -6069
rect 53250 -6121 53260 -6069
rect 53380 -6121 53390 -6069
rect 53442 -6121 53452 -6069
rect 53571 -6122 53581 -6070
rect 53633 -6122 53643 -6070
rect 53766 -6122 53776 -6070
rect 53828 -6122 53838 -6070
rect 53956 -6122 53966 -6070
rect 54018 -6122 54028 -6070
rect 54147 -6122 54157 -6070
rect 54209 -6122 54219 -6070
rect 54339 -6122 54349 -6070
rect 54401 -6122 54411 -6070
rect 54532 -6121 54542 -6069
rect 54594 -6121 54604 -6069
rect 54724 -6122 54734 -6070
rect 54786 -6122 54796 -6070
rect 54916 -6122 54926 -6070
rect 54978 -6122 54988 -6070
rect 55109 -6122 55119 -6070
rect 55171 -6122 55181 -6070
rect 55300 -6121 55310 -6069
rect 55362 -6121 55372 -6069
rect 55492 -6122 55502 -6070
rect 55554 -6122 55564 -6070
rect 55684 -6121 55694 -6069
rect 55746 -6121 55756 -6069
rect 55876 -6121 55886 -6069
rect 55938 -6121 55948 -6069
rect 56067 -6122 56077 -6070
rect 56129 -6122 56139 -6070
rect 56260 -6121 56270 -6069
rect 56322 -6121 56332 -6069
rect 56452 -6121 56462 -6069
rect 56514 -6121 56524 -6069
rect 56646 -6122 56656 -6070
rect 56708 -6122 56718 -6070
rect 56837 -6123 56847 -6071
rect 56899 -6123 56909 -6071
rect 57026 -6122 57036 -6070
rect 57088 -6122 57098 -6070
rect 57219 -6122 57229 -6070
rect 57281 -6122 57291 -6070
rect 57412 -6122 57422 -6070
rect 57474 -6122 57484 -6070
rect 57603 -6121 57613 -6069
rect 57665 -6121 57675 -6069
rect 57794 -6121 57804 -6069
rect 57856 -6121 57866 -6069
rect 51939 -6262 51949 -6210
rect 52001 -6262 52011 -6210
rect 52131 -6262 52141 -6210
rect 52193 -6262 52203 -6210
rect 52324 -6262 52334 -6210
rect 52386 -6262 52396 -6210
rect 52516 -6262 52526 -6210
rect 52578 -6262 52588 -6210
rect 52709 -6262 52719 -6210
rect 52771 -6262 52781 -6210
rect 52901 -6261 52911 -6209
rect 52963 -6261 52973 -6209
rect 53092 -6262 53102 -6210
rect 53154 -6262 53164 -6210
rect 53284 -6262 53294 -6210
rect 53346 -6262 53356 -6210
rect 53476 -6261 53486 -6209
rect 53538 -6261 53548 -6209
rect 53668 -6261 53678 -6209
rect 53730 -6261 53740 -6209
rect 53860 -6262 53870 -6210
rect 53922 -6262 53932 -6210
rect 54052 -6261 54062 -6209
rect 54114 -6261 54124 -6209
rect 54244 -6262 54254 -6210
rect 54306 -6262 54316 -6210
rect 54435 -6261 54445 -6209
rect 54497 -6261 54507 -6209
rect 54629 -6262 54639 -6210
rect 54691 -6262 54701 -6210
rect 54819 -6262 54829 -6210
rect 54881 -6262 54891 -6210
rect 55011 -6262 55021 -6210
rect 55073 -6262 55083 -6210
rect 55204 -6262 55214 -6210
rect 55266 -6262 55276 -6210
rect 55395 -6262 55405 -6210
rect 55457 -6262 55467 -6210
rect 55588 -6261 55598 -6209
rect 55650 -6261 55660 -6209
rect 55781 -6262 55791 -6210
rect 55843 -6262 55853 -6210
rect 55972 -6262 55982 -6210
rect 56034 -6262 56044 -6210
rect 56165 -6262 56175 -6210
rect 56227 -6262 56237 -6210
rect 56355 -6262 56365 -6210
rect 56417 -6262 56427 -6210
rect 56549 -6261 56559 -6209
rect 56611 -6261 56621 -6209
rect 56738 -6262 56748 -6210
rect 56800 -6262 56810 -6210
rect 56931 -6262 56941 -6210
rect 56993 -6262 57003 -6210
rect 57124 -6262 57134 -6210
rect 57186 -6262 57196 -6210
rect 57314 -6262 57324 -6210
rect 57376 -6262 57386 -6210
rect 57507 -6261 57517 -6209
rect 57569 -6261 57579 -6209
rect 57696 -6261 57706 -6209
rect 57758 -6261 57768 -6209
rect 57910 -6300 57940 -6020
rect 51860 -6310 57940 -6300
rect 51860 -6320 57800 -6310
rect 50970 -6368 51328 -6326
rect 51860 -6330 52040 -6320
rect 50970 -6456 51016 -6368
rect 51106 -6448 51116 -6396
rect 51168 -6448 51178 -6396
rect 51286 -6446 51328 -6368
rect 52030 -6380 52040 -6330
rect 52100 -6330 57800 -6320
rect 52100 -6380 52110 -6330
rect 57790 -6370 57800 -6330
rect 57860 -6330 57940 -6310
rect 58070 -6020 64130 -5990
rect 66908 -6002 66918 -5950
rect 66970 -6002 66980 -5950
rect 58070 -6300 58100 -6020
rect 58231 -6122 58241 -6070
rect 58293 -6122 58303 -6070
rect 58421 -6121 58431 -6069
rect 58483 -6121 58493 -6069
rect 58613 -6120 58623 -6068
rect 58675 -6120 58685 -6068
rect 58804 -6120 58814 -6068
rect 58866 -6120 58876 -6068
rect 58998 -6120 59008 -6068
rect 59060 -6120 59070 -6068
rect 59188 -6121 59198 -6069
rect 59250 -6121 59260 -6069
rect 59382 -6120 59392 -6068
rect 59444 -6120 59454 -6068
rect 59574 -6120 59584 -6068
rect 59636 -6120 59646 -6068
rect 59765 -6121 59775 -6069
rect 59827 -6121 59837 -6069
rect 59960 -6121 59970 -6069
rect 60022 -6121 60032 -6069
rect 60150 -6121 60160 -6069
rect 60212 -6121 60222 -6069
rect 60341 -6121 60351 -6069
rect 60403 -6121 60413 -6069
rect 60533 -6121 60543 -6069
rect 60595 -6121 60605 -6069
rect 60726 -6120 60736 -6068
rect 60788 -6120 60798 -6068
rect 60918 -6121 60928 -6069
rect 60980 -6121 60990 -6069
rect 61110 -6121 61120 -6069
rect 61172 -6121 61182 -6069
rect 61303 -6121 61313 -6069
rect 61365 -6121 61375 -6069
rect 61494 -6120 61504 -6068
rect 61556 -6120 61566 -6068
rect 61686 -6121 61696 -6069
rect 61748 -6121 61758 -6069
rect 61878 -6120 61888 -6068
rect 61940 -6120 61950 -6068
rect 62070 -6120 62080 -6068
rect 62132 -6120 62142 -6068
rect 62261 -6121 62271 -6069
rect 62323 -6121 62333 -6069
rect 62454 -6120 62464 -6068
rect 62516 -6120 62526 -6068
rect 62646 -6120 62656 -6068
rect 62708 -6120 62718 -6068
rect 62840 -6121 62850 -6069
rect 62902 -6121 62912 -6069
rect 63031 -6122 63041 -6070
rect 63093 -6122 63103 -6070
rect 63220 -6121 63230 -6069
rect 63282 -6121 63292 -6069
rect 63413 -6121 63423 -6069
rect 63475 -6121 63485 -6069
rect 63606 -6121 63616 -6069
rect 63668 -6121 63678 -6069
rect 63797 -6120 63807 -6068
rect 63859 -6120 63869 -6068
rect 63988 -6120 63998 -6068
rect 64050 -6120 64060 -6068
rect 58133 -6261 58143 -6209
rect 58195 -6261 58205 -6209
rect 58325 -6261 58335 -6209
rect 58387 -6261 58397 -6209
rect 58518 -6261 58528 -6209
rect 58580 -6261 58590 -6209
rect 58710 -6261 58720 -6209
rect 58772 -6261 58782 -6209
rect 58903 -6261 58913 -6209
rect 58965 -6261 58975 -6209
rect 59095 -6260 59105 -6208
rect 59157 -6260 59167 -6208
rect 59286 -6261 59296 -6209
rect 59348 -6261 59358 -6209
rect 59478 -6261 59488 -6209
rect 59540 -6261 59550 -6209
rect 59670 -6260 59680 -6208
rect 59732 -6260 59742 -6208
rect 59862 -6260 59872 -6208
rect 59924 -6260 59934 -6208
rect 60054 -6261 60064 -6209
rect 60116 -6261 60126 -6209
rect 60246 -6260 60256 -6208
rect 60308 -6260 60318 -6208
rect 60438 -6261 60448 -6209
rect 60500 -6261 60510 -6209
rect 60629 -6260 60639 -6208
rect 60691 -6260 60701 -6208
rect 60823 -6261 60833 -6209
rect 60885 -6261 60895 -6209
rect 61013 -6261 61023 -6209
rect 61075 -6261 61085 -6209
rect 61205 -6261 61215 -6209
rect 61267 -6261 61277 -6209
rect 61398 -6261 61408 -6209
rect 61460 -6261 61470 -6209
rect 61589 -6261 61599 -6209
rect 61651 -6261 61661 -6209
rect 61782 -6260 61792 -6208
rect 61844 -6260 61854 -6208
rect 61975 -6261 61985 -6209
rect 62037 -6261 62047 -6209
rect 62166 -6261 62176 -6209
rect 62228 -6261 62238 -6209
rect 62359 -6261 62369 -6209
rect 62421 -6261 62431 -6209
rect 62549 -6261 62559 -6209
rect 62611 -6261 62621 -6209
rect 62743 -6260 62753 -6208
rect 62805 -6260 62815 -6208
rect 62932 -6261 62942 -6209
rect 62994 -6261 63004 -6209
rect 63125 -6261 63135 -6209
rect 63187 -6261 63197 -6209
rect 63318 -6261 63328 -6209
rect 63380 -6261 63390 -6209
rect 63508 -6261 63518 -6209
rect 63570 -6261 63580 -6209
rect 63701 -6260 63711 -6208
rect 63763 -6260 63773 -6208
rect 63890 -6260 63900 -6208
rect 63952 -6260 63962 -6208
rect 64100 -6300 64130 -6020
rect 68000 -6298 68362 -5710
rect 68920 -6272 68930 -5188
rect 69296 -6272 69306 -5188
rect 58070 -6310 63990 -6300
rect 58070 -6330 58230 -6310
rect 57860 -6370 57870 -6330
rect 58220 -6370 58230 -6330
rect 58290 -6330 63990 -6310
rect 58290 -6370 58300 -6330
rect 63980 -6360 63990 -6330
rect 64050 -6330 64130 -6300
rect 64050 -6360 64060 -6330
rect 64382 -6340 64738 -6302
rect 64382 -6446 64424 -6340
rect 64520 -6432 64530 -6380
rect 64582 -6432 64592 -6380
rect 51286 -6490 64424 -6446
rect 64690 -6458 64736 -6340
rect 51106 -6552 51116 -6500
rect 51168 -6552 51178 -6500
rect 64526 -6548 64536 -6496
rect 64588 -6548 64598 -6496
rect 51874 -6640 57930 -6610
rect 47244 -7752 47254 -6678
rect 47614 -7752 47624 -6678
rect 48194 -7240 48556 -6644
rect 49426 -6924 49436 -6872
rect 49488 -6924 49498 -6872
rect 51874 -6920 51904 -6640
rect 52038 -6741 52048 -6689
rect 52100 -6741 52110 -6689
rect 52228 -6740 52238 -6688
rect 52290 -6740 52300 -6688
rect 52420 -6739 52430 -6687
rect 52482 -6739 52492 -6687
rect 52611 -6739 52621 -6687
rect 52673 -6739 52683 -6687
rect 52805 -6739 52815 -6687
rect 52867 -6739 52877 -6687
rect 52995 -6740 53005 -6688
rect 53057 -6740 53067 -6688
rect 53189 -6739 53199 -6687
rect 53251 -6739 53261 -6687
rect 53381 -6739 53391 -6687
rect 53443 -6739 53453 -6687
rect 53572 -6740 53582 -6688
rect 53634 -6740 53644 -6688
rect 53767 -6740 53777 -6688
rect 53829 -6740 53839 -6688
rect 53957 -6740 53967 -6688
rect 54019 -6740 54029 -6688
rect 54148 -6740 54158 -6688
rect 54210 -6740 54220 -6688
rect 54340 -6740 54350 -6688
rect 54402 -6740 54412 -6688
rect 54533 -6739 54543 -6687
rect 54595 -6739 54605 -6687
rect 54725 -6740 54735 -6688
rect 54787 -6740 54797 -6688
rect 54917 -6740 54927 -6688
rect 54979 -6740 54989 -6688
rect 55110 -6740 55120 -6688
rect 55172 -6740 55182 -6688
rect 55301 -6739 55311 -6687
rect 55363 -6739 55373 -6687
rect 55493 -6740 55503 -6688
rect 55555 -6740 55565 -6688
rect 55685 -6739 55695 -6687
rect 55747 -6739 55757 -6687
rect 55877 -6739 55887 -6687
rect 55939 -6739 55949 -6687
rect 56068 -6740 56078 -6688
rect 56130 -6740 56140 -6688
rect 56261 -6739 56271 -6687
rect 56323 -6739 56333 -6687
rect 56453 -6739 56463 -6687
rect 56515 -6739 56525 -6687
rect 56647 -6740 56657 -6688
rect 56709 -6740 56719 -6688
rect 56838 -6741 56848 -6689
rect 56900 -6741 56910 -6689
rect 57027 -6740 57037 -6688
rect 57089 -6740 57099 -6688
rect 57220 -6740 57230 -6688
rect 57282 -6740 57292 -6688
rect 57413 -6740 57423 -6688
rect 57475 -6740 57485 -6688
rect 57604 -6739 57614 -6687
rect 57666 -6739 57676 -6687
rect 57795 -6739 57805 -6687
rect 57857 -6739 57867 -6687
rect 51940 -6880 51950 -6828
rect 52002 -6880 52012 -6828
rect 52132 -6880 52142 -6828
rect 52194 -6880 52204 -6828
rect 52325 -6880 52335 -6828
rect 52387 -6880 52397 -6828
rect 52517 -6880 52527 -6828
rect 52579 -6880 52589 -6828
rect 52710 -6880 52720 -6828
rect 52772 -6880 52782 -6828
rect 52902 -6879 52912 -6827
rect 52964 -6879 52974 -6827
rect 53093 -6880 53103 -6828
rect 53155 -6880 53165 -6828
rect 53285 -6880 53295 -6828
rect 53347 -6880 53357 -6828
rect 53477 -6879 53487 -6827
rect 53539 -6879 53549 -6827
rect 53669 -6879 53679 -6827
rect 53731 -6879 53741 -6827
rect 53861 -6880 53871 -6828
rect 53923 -6880 53933 -6828
rect 54053 -6879 54063 -6827
rect 54115 -6879 54125 -6827
rect 54245 -6880 54255 -6828
rect 54307 -6880 54317 -6828
rect 54436 -6879 54446 -6827
rect 54498 -6879 54508 -6827
rect 54630 -6880 54640 -6828
rect 54692 -6880 54702 -6828
rect 54820 -6880 54830 -6828
rect 54882 -6880 54892 -6828
rect 55012 -6880 55022 -6828
rect 55074 -6880 55084 -6828
rect 55205 -6880 55215 -6828
rect 55267 -6880 55277 -6828
rect 55396 -6880 55406 -6828
rect 55458 -6880 55468 -6828
rect 55589 -6879 55599 -6827
rect 55651 -6879 55661 -6827
rect 55782 -6880 55792 -6828
rect 55844 -6880 55854 -6828
rect 55973 -6880 55983 -6828
rect 56035 -6880 56045 -6828
rect 56166 -6880 56176 -6828
rect 56228 -6880 56238 -6828
rect 56356 -6880 56366 -6828
rect 56418 -6880 56428 -6828
rect 56550 -6879 56560 -6827
rect 56612 -6879 56622 -6827
rect 56739 -6880 56749 -6828
rect 56801 -6880 56811 -6828
rect 56932 -6880 56942 -6828
rect 56994 -6880 57004 -6828
rect 57125 -6880 57135 -6828
rect 57187 -6880 57197 -6828
rect 57315 -6880 57325 -6828
rect 57377 -6880 57387 -6828
rect 57508 -6879 57518 -6827
rect 57570 -6879 57580 -6827
rect 57697 -6879 57707 -6827
rect 57759 -6879 57769 -6827
rect 57900 -6920 57930 -6640
rect 51874 -6950 57930 -6920
rect 58070 -6640 64114 -6610
rect 58070 -6920 58100 -6640
rect 58226 -6740 58236 -6688
rect 58288 -6740 58298 -6688
rect 58416 -6739 58426 -6687
rect 58478 -6739 58488 -6687
rect 58608 -6738 58618 -6686
rect 58670 -6738 58680 -6686
rect 58799 -6738 58809 -6686
rect 58861 -6738 58871 -6686
rect 58993 -6738 59003 -6686
rect 59055 -6738 59065 -6686
rect 59183 -6739 59193 -6687
rect 59245 -6739 59255 -6687
rect 59377 -6738 59387 -6686
rect 59439 -6738 59449 -6686
rect 59569 -6738 59579 -6686
rect 59631 -6738 59641 -6686
rect 59760 -6739 59770 -6687
rect 59822 -6739 59832 -6687
rect 59955 -6739 59965 -6687
rect 60017 -6739 60027 -6687
rect 60145 -6739 60155 -6687
rect 60207 -6739 60217 -6687
rect 60336 -6739 60346 -6687
rect 60398 -6739 60408 -6687
rect 60528 -6739 60538 -6687
rect 60590 -6739 60600 -6687
rect 60721 -6738 60731 -6686
rect 60783 -6738 60793 -6686
rect 60913 -6739 60923 -6687
rect 60975 -6739 60985 -6687
rect 61105 -6739 61115 -6687
rect 61167 -6739 61177 -6687
rect 61298 -6739 61308 -6687
rect 61360 -6739 61370 -6687
rect 61489 -6738 61499 -6686
rect 61551 -6738 61561 -6686
rect 61681 -6739 61691 -6687
rect 61743 -6739 61753 -6687
rect 61873 -6738 61883 -6686
rect 61935 -6738 61945 -6686
rect 62065 -6738 62075 -6686
rect 62127 -6738 62137 -6686
rect 62256 -6739 62266 -6687
rect 62318 -6739 62328 -6687
rect 62449 -6738 62459 -6686
rect 62511 -6738 62521 -6686
rect 62641 -6738 62651 -6686
rect 62703 -6738 62713 -6686
rect 62835 -6739 62845 -6687
rect 62897 -6739 62907 -6687
rect 63026 -6740 63036 -6688
rect 63088 -6740 63098 -6688
rect 63215 -6739 63225 -6687
rect 63277 -6739 63287 -6687
rect 63408 -6739 63418 -6687
rect 63470 -6739 63480 -6687
rect 63601 -6739 63611 -6687
rect 63663 -6739 63673 -6687
rect 63792 -6738 63802 -6686
rect 63854 -6738 63864 -6686
rect 63983 -6738 63993 -6686
rect 64045 -6738 64055 -6686
rect 58130 -6879 58138 -6827
rect 58190 -6879 58200 -6827
rect 58320 -6879 58330 -6827
rect 58382 -6879 58392 -6827
rect 58513 -6879 58523 -6827
rect 58575 -6879 58585 -6827
rect 58705 -6879 58715 -6827
rect 58767 -6879 58777 -6827
rect 58898 -6879 58908 -6827
rect 58960 -6879 58970 -6827
rect 59090 -6878 59100 -6826
rect 59152 -6878 59162 -6826
rect 59281 -6879 59291 -6827
rect 59343 -6879 59353 -6827
rect 59473 -6879 59483 -6827
rect 59535 -6879 59545 -6827
rect 59665 -6878 59675 -6826
rect 59727 -6878 59737 -6826
rect 59857 -6878 59867 -6826
rect 59919 -6878 59929 -6826
rect 60049 -6879 60059 -6827
rect 60111 -6879 60121 -6827
rect 60241 -6878 60251 -6826
rect 60303 -6878 60313 -6826
rect 60433 -6879 60443 -6827
rect 60495 -6879 60505 -6827
rect 60624 -6878 60634 -6826
rect 60686 -6878 60696 -6826
rect 60818 -6879 60828 -6827
rect 60880 -6879 60890 -6827
rect 61008 -6879 61018 -6827
rect 61070 -6879 61080 -6827
rect 61200 -6879 61210 -6827
rect 61262 -6879 61272 -6827
rect 61393 -6879 61403 -6827
rect 61455 -6879 61465 -6827
rect 61584 -6879 61594 -6827
rect 61646 -6879 61656 -6827
rect 61777 -6878 61787 -6826
rect 61839 -6878 61849 -6826
rect 61970 -6879 61980 -6827
rect 62032 -6879 62042 -6827
rect 62161 -6879 62171 -6827
rect 62223 -6879 62233 -6827
rect 62354 -6879 62364 -6827
rect 62416 -6879 62426 -6827
rect 62544 -6879 62554 -6827
rect 62606 -6879 62616 -6827
rect 62738 -6878 62748 -6826
rect 62800 -6878 62810 -6826
rect 62927 -6879 62937 -6827
rect 62989 -6879 62999 -6827
rect 63120 -6879 63130 -6827
rect 63182 -6879 63192 -6827
rect 63313 -6879 63323 -6827
rect 63375 -6879 63385 -6827
rect 63503 -6879 63513 -6827
rect 63565 -6879 63575 -6827
rect 63696 -6878 63706 -6826
rect 63758 -6878 63768 -6826
rect 63885 -6878 63895 -6826
rect 63947 -6878 63957 -6826
rect 64084 -6920 64114 -6640
rect 66902 -6902 66912 -6850
rect 66964 -6902 66974 -6850
rect 58070 -6950 64114 -6920
rect 48190 -7640 48556 -7240
rect 49890 -7260 66624 -7230
rect 49890 -7540 49920 -7260
rect 50077 -7354 50087 -7302
rect 50139 -7354 50149 -7302
rect 50267 -7353 50277 -7301
rect 50329 -7353 50339 -7301
rect 50460 -7356 50470 -7304
rect 50522 -7356 50532 -7304
rect 50652 -7351 50662 -7299
rect 50714 -7351 50724 -7299
rect 50844 -7355 50854 -7303
rect 50906 -7355 50916 -7303
rect 51036 -7350 51046 -7298
rect 51098 -7350 51108 -7298
rect 51228 -7351 51238 -7299
rect 51290 -7351 51300 -7299
rect 51418 -7350 51428 -7298
rect 51480 -7350 51490 -7298
rect 51612 -7361 51622 -7309
rect 51674 -7361 51684 -7309
rect 51801 -7359 51811 -7307
rect 51863 -7359 51873 -7307
rect 51991 -7359 52001 -7307
rect 52053 -7359 52063 -7307
rect 52190 -7360 52200 -7308
rect 52252 -7360 52262 -7308
rect 52382 -7359 52392 -7307
rect 52444 -7359 52454 -7307
rect 52572 -7360 52582 -7308
rect 52634 -7360 52644 -7308
rect 52764 -7353 52774 -7301
rect 52826 -7353 52836 -7301
rect 52956 -7303 53028 -7298
rect 52956 -7355 52966 -7303
rect 53018 -7355 53028 -7303
rect 53149 -7354 53159 -7302
rect 53211 -7354 53221 -7302
rect 53341 -7352 53351 -7300
rect 53403 -7352 53413 -7300
rect 53532 -7352 53542 -7300
rect 53594 -7352 53604 -7300
rect 53726 -7357 53736 -7305
rect 53788 -7357 53798 -7305
rect 53917 -7353 53927 -7301
rect 53979 -7353 53989 -7301
rect 54109 -7349 54119 -7297
rect 54171 -7349 54181 -7297
rect 54302 -7353 54312 -7301
rect 54364 -7353 54374 -7301
rect 54494 -7353 54504 -7301
rect 54556 -7353 54566 -7301
rect 54687 -7354 54697 -7302
rect 54749 -7354 54759 -7302
rect 54879 -7352 54889 -7300
rect 54941 -7352 54951 -7300
rect 55070 -7351 55080 -7299
rect 55132 -7351 55142 -7299
rect 55261 -7350 55271 -7298
rect 55323 -7350 55333 -7298
rect 55454 -7350 55464 -7298
rect 55516 -7350 55526 -7298
rect 55645 -7359 55655 -7307
rect 55707 -7359 55717 -7307
rect 55836 -7360 55846 -7308
rect 55898 -7360 55908 -7308
rect 56026 -7361 56036 -7309
rect 56088 -7361 56098 -7309
rect 56220 -7365 56230 -7313
rect 56282 -7365 56292 -7313
rect 56412 -7367 56422 -7315
rect 56474 -7367 56484 -7315
rect 56606 -7366 56616 -7314
rect 56668 -7366 56678 -7314
rect 56798 -7363 56808 -7311
rect 56860 -7363 56870 -7311
rect 56987 -7360 56997 -7308
rect 57049 -7360 57059 -7308
rect 57181 -7358 57191 -7306
rect 57243 -7358 57253 -7306
rect 57374 -7359 57384 -7307
rect 57436 -7359 57446 -7307
rect 57567 -7360 57577 -7308
rect 57629 -7360 57639 -7308
rect 57756 -7360 57766 -7308
rect 57818 -7360 57828 -7308
rect 57949 -7360 57959 -7308
rect 58011 -7360 58021 -7308
rect 58141 -7360 58151 -7308
rect 58203 -7360 58213 -7308
rect 58332 -7360 58342 -7308
rect 58394 -7360 58404 -7308
rect 58525 -7360 58535 -7308
rect 58587 -7360 58597 -7308
rect 58716 -7359 58726 -7307
rect 58778 -7359 58788 -7307
rect 58911 -7360 58921 -7308
rect 58973 -7360 58983 -7308
rect 59100 -7360 59110 -7308
rect 59162 -7360 59172 -7308
rect 59293 -7360 59303 -7308
rect 59355 -7360 59365 -7308
rect 59485 -7360 59495 -7308
rect 59547 -7360 59557 -7308
rect 59676 -7360 59686 -7308
rect 59738 -7360 59748 -7308
rect 59868 -7360 59878 -7308
rect 59930 -7360 59940 -7308
rect 60061 -7360 60071 -7308
rect 60123 -7360 60133 -7308
rect 60250 -7361 60260 -7309
rect 60312 -7361 60322 -7309
rect 60444 -7360 60454 -7308
rect 60506 -7360 60516 -7308
rect 60635 -7360 60645 -7308
rect 60697 -7360 60707 -7308
rect 60828 -7360 60838 -7308
rect 60890 -7360 60900 -7308
rect 61020 -7360 61030 -7308
rect 61082 -7360 61092 -7308
rect 61212 -7361 61222 -7309
rect 61274 -7361 61284 -7309
rect 61405 -7359 61415 -7307
rect 61467 -7359 61477 -7307
rect 61595 -7359 61605 -7307
rect 61657 -7359 61667 -7307
rect 61788 -7361 61798 -7309
rect 61850 -7361 61860 -7309
rect 61980 -7360 61990 -7308
rect 62042 -7360 62052 -7308
rect 62173 -7359 62183 -7307
rect 62235 -7359 62245 -7307
rect 62364 -7359 62374 -7307
rect 62426 -7359 62436 -7307
rect 62556 -7360 62566 -7308
rect 62618 -7360 62628 -7308
rect 62747 -7360 62757 -7308
rect 62809 -7360 62819 -7308
rect 62939 -7360 62949 -7308
rect 63001 -7360 63011 -7308
rect 63133 -7359 63143 -7307
rect 63195 -7359 63205 -7307
rect 63325 -7360 63335 -7308
rect 63387 -7360 63397 -7308
rect 63515 -7361 63525 -7309
rect 63577 -7361 63587 -7309
rect 63706 -7362 63716 -7310
rect 63768 -7362 63778 -7310
rect 63899 -7360 63909 -7308
rect 63961 -7360 63971 -7308
rect 64092 -7359 64102 -7307
rect 64154 -7359 64164 -7307
rect 64285 -7360 64295 -7308
rect 64347 -7360 64357 -7308
rect 64476 -7360 64486 -7308
rect 64538 -7360 64548 -7308
rect 64667 -7360 64677 -7308
rect 64729 -7360 64739 -7308
rect 64860 -7360 64870 -7308
rect 64922 -7360 64932 -7308
rect 65053 -7360 65063 -7308
rect 65115 -7360 65125 -7308
rect 65244 -7360 65254 -7308
rect 65306 -7360 65316 -7308
rect 65435 -7359 65445 -7307
rect 65497 -7359 65507 -7307
rect 65626 -7359 65636 -7307
rect 65688 -7359 65698 -7307
rect 65819 -7360 65829 -7308
rect 65881 -7360 65891 -7308
rect 66013 -7360 66023 -7308
rect 66075 -7360 66085 -7308
rect 66201 -7361 66211 -7309
rect 66263 -7361 66273 -7309
rect 66395 -7369 66405 -7317
rect 66457 -7369 66467 -7317
rect 49981 -7497 49991 -7445
rect 50043 -7497 50053 -7445
rect 50172 -7499 50182 -7447
rect 50234 -7499 50244 -7447
rect 50364 -7498 50374 -7446
rect 50426 -7498 50436 -7446
rect 50556 -7501 50566 -7449
rect 50618 -7501 50628 -7449
rect 50750 -7500 50760 -7448
rect 50812 -7500 50822 -7448
rect 50940 -7500 50950 -7448
rect 51002 -7500 51012 -7448
rect 51135 -7498 51145 -7446
rect 51197 -7498 51207 -7446
rect 51326 -7497 51336 -7445
rect 51388 -7497 51398 -7445
rect 51521 -7499 51531 -7447
rect 51583 -7499 51593 -7447
rect 51711 -7499 51721 -7447
rect 51773 -7499 51783 -7447
rect 51901 -7498 51911 -7446
rect 51963 -7498 51973 -7446
rect 52094 -7497 52104 -7445
rect 52156 -7497 52166 -7445
rect 52285 -7497 52295 -7445
rect 52347 -7497 52357 -7445
rect 52481 -7499 52491 -7447
rect 52543 -7499 52553 -7447
rect 52670 -7499 52680 -7447
rect 52732 -7499 52742 -7447
rect 52864 -7499 52874 -7447
rect 52926 -7499 52936 -7447
rect 53053 -7499 53063 -7447
rect 53115 -7499 53125 -7447
rect 53245 -7500 53255 -7448
rect 53307 -7500 53317 -7448
rect 53438 -7500 53448 -7448
rect 53500 -7500 53510 -7448
rect 53629 -7500 53639 -7448
rect 53691 -7500 53701 -7448
rect 53821 -7499 53831 -7447
rect 53883 -7499 53893 -7447
rect 54013 -7500 54023 -7448
rect 54075 -7500 54085 -7448
rect 54206 -7500 54216 -7448
rect 54268 -7500 54278 -7448
rect 54397 -7500 54407 -7448
rect 54459 -7500 54469 -7448
rect 54589 -7499 54599 -7447
rect 54651 -7499 54661 -7447
rect 54782 -7500 54792 -7448
rect 54844 -7500 54854 -7448
rect 54974 -7500 54984 -7448
rect 55036 -7500 55046 -7448
rect 55165 -7500 55175 -7448
rect 55227 -7500 55237 -7448
rect 55356 -7500 55366 -7448
rect 55418 -7500 55428 -7448
rect 55548 -7500 55558 -7448
rect 55610 -7500 55620 -7448
rect 55741 -7499 55751 -7447
rect 55803 -7499 55813 -7447
rect 55932 -7499 55942 -7447
rect 55994 -7499 56004 -7447
rect 56126 -7500 56136 -7448
rect 56188 -7500 56198 -7448
rect 56318 -7500 56328 -7448
rect 56380 -7500 56390 -7448
rect 56510 -7500 56520 -7448
rect 56572 -7500 56582 -7448
rect 56702 -7500 56712 -7448
rect 56764 -7500 56774 -7448
rect 56894 -7500 56904 -7448
rect 56956 -7500 56966 -7448
rect 57086 -7500 57096 -7448
rect 57148 -7500 57158 -7448
rect 57278 -7500 57288 -7448
rect 57340 -7500 57350 -7448
rect 57469 -7500 57479 -7448
rect 57531 -7500 57541 -7448
rect 57661 -7500 57671 -7448
rect 57723 -7500 57733 -7448
rect 57854 -7500 57864 -7448
rect 57916 -7500 57926 -7448
rect 58046 -7500 58056 -7448
rect 58108 -7500 58118 -7448
rect 58238 -7500 58248 -7448
rect 58300 -7500 58310 -7448
rect 58429 -7500 58439 -7448
rect 58491 -7500 58501 -7448
rect 58621 -7500 58631 -7448
rect 58683 -7500 58693 -7448
rect 58812 -7500 58822 -7448
rect 58874 -7500 58884 -7448
rect 59003 -7500 59013 -7448
rect 59065 -7500 59075 -7448
rect 59197 -7500 59207 -7448
rect 59259 -7500 59269 -7448
rect 59389 -7500 59399 -7448
rect 59451 -7500 59461 -7448
rect 59582 -7499 59592 -7447
rect 59644 -7499 59654 -7447
rect 59773 -7500 59783 -7448
rect 59835 -7500 59845 -7448
rect 59965 -7500 59975 -7448
rect 60027 -7500 60037 -7448
rect 60158 -7500 60168 -7448
rect 60220 -7500 60230 -7448
rect 60350 -7500 60360 -7448
rect 60412 -7500 60422 -7448
rect 60543 -7499 60553 -7447
rect 60605 -7499 60615 -7447
rect 60734 -7500 60744 -7448
rect 60796 -7500 60806 -7448
rect 60926 -7500 60936 -7448
rect 60988 -7500 60998 -7448
rect 61117 -7500 61127 -7448
rect 61179 -7500 61189 -7448
rect 61309 -7500 61319 -7448
rect 61371 -7500 61381 -7448
rect 61501 -7500 61511 -7448
rect 61563 -7500 61573 -7448
rect 61694 -7500 61704 -7448
rect 61756 -7500 61766 -7448
rect 61885 -7500 61895 -7448
rect 61947 -7500 61957 -7448
rect 62077 -7500 62087 -7448
rect 62139 -7500 62149 -7448
rect 62269 -7499 62279 -7447
rect 62331 -7499 62341 -7447
rect 62461 -7500 62471 -7448
rect 62523 -7500 62533 -7448
rect 62651 -7500 62661 -7448
rect 62713 -7500 62723 -7448
rect 62845 -7500 62855 -7448
rect 62907 -7500 62917 -7448
rect 63037 -7499 63047 -7447
rect 63099 -7499 63109 -7447
rect 63228 -7500 63238 -7448
rect 63290 -7500 63300 -7448
rect 63421 -7500 63431 -7448
rect 63483 -7500 63493 -7448
rect 63612 -7499 63622 -7447
rect 63674 -7499 63684 -7447
rect 63804 -7500 63814 -7448
rect 63866 -7500 63876 -7448
rect 63995 -7500 64005 -7448
rect 64057 -7500 64067 -7448
rect 64189 -7499 64199 -7447
rect 64251 -7499 64261 -7447
rect 64380 -7500 64390 -7448
rect 64442 -7500 64452 -7448
rect 64572 -7500 64582 -7448
rect 64634 -7500 64644 -7448
rect 64764 -7500 64774 -7448
rect 64826 -7500 64836 -7448
rect 64956 -7500 64966 -7448
rect 65018 -7500 65028 -7448
rect 65149 -7500 65159 -7448
rect 65211 -7500 65221 -7448
rect 65340 -7500 65350 -7448
rect 65402 -7500 65412 -7448
rect 65533 -7499 65543 -7447
rect 65595 -7499 65605 -7447
rect 65724 -7500 65734 -7448
rect 65786 -7500 65796 -7448
rect 65917 -7500 65927 -7448
rect 65979 -7500 65989 -7448
rect 66108 -7500 66118 -7448
rect 66170 -7500 66180 -7448
rect 66299 -7498 66309 -7446
rect 66361 -7498 66371 -7446
rect 66494 -7500 66504 -7448
rect 66556 -7500 66566 -7448
rect 66594 -7540 66624 -7260
rect 49890 -7570 66624 -7540
rect 68006 -7234 68368 -6644
rect 68006 -7640 68374 -7234
rect 68368 -7642 68374 -7640
rect 49928 -7664 66600 -7658
rect 48262 -7706 48458 -7700
rect 48262 -7764 48274 -7706
rect 48446 -7764 48458 -7706
rect 49928 -7756 49940 -7664
rect 66588 -7756 66600 -7664
rect 49928 -7762 66600 -7756
rect 68108 -7710 68304 -7704
rect 48262 -7770 48458 -7764
rect 68108 -7768 68120 -7710
rect 68292 -7768 68304 -7710
rect 68914 -7756 68924 -6672
rect 69290 -7756 69300 -6672
rect 68108 -7774 68304 -7768
<< via1 >>
rect 47260 -6264 47620 -5190
rect 48286 -5236 48458 -5178
rect 49920 -5280 66568 -5188
rect 68070 -5236 68242 -5178
rect 50087 -5494 50139 -5442
rect 50277 -5493 50329 -5441
rect 50470 -5496 50522 -5444
rect 50662 -5491 50714 -5439
rect 50854 -5495 50906 -5443
rect 51046 -5490 51098 -5438
rect 51238 -5491 51290 -5439
rect 51428 -5490 51480 -5438
rect 51622 -5501 51674 -5449
rect 51811 -5499 51863 -5447
rect 52001 -5499 52053 -5447
rect 52200 -5500 52252 -5448
rect 52392 -5499 52444 -5447
rect 52582 -5500 52634 -5448
rect 52774 -5493 52826 -5441
rect 52966 -5495 53018 -5443
rect 53159 -5494 53211 -5442
rect 53351 -5492 53403 -5440
rect 53542 -5492 53594 -5440
rect 53736 -5497 53788 -5445
rect 53927 -5493 53979 -5441
rect 54119 -5489 54171 -5437
rect 54312 -5493 54364 -5441
rect 54504 -5493 54556 -5441
rect 54697 -5494 54749 -5442
rect 54889 -5492 54941 -5440
rect 55080 -5491 55132 -5439
rect 55271 -5490 55323 -5438
rect 55464 -5490 55516 -5438
rect 55655 -5499 55707 -5447
rect 55846 -5500 55898 -5448
rect 56036 -5501 56088 -5449
rect 56230 -5505 56282 -5453
rect 56422 -5507 56474 -5455
rect 56616 -5506 56668 -5454
rect 56808 -5503 56860 -5451
rect 56997 -5500 57049 -5448
rect 57191 -5498 57243 -5446
rect 57384 -5499 57436 -5447
rect 57577 -5500 57629 -5448
rect 57766 -5500 57818 -5448
rect 57959 -5500 58011 -5448
rect 58151 -5500 58203 -5448
rect 58342 -5500 58394 -5448
rect 58535 -5500 58587 -5448
rect 58726 -5499 58778 -5447
rect 58921 -5500 58973 -5448
rect 59110 -5500 59162 -5448
rect 59303 -5500 59355 -5448
rect 59495 -5500 59547 -5448
rect 59686 -5500 59738 -5448
rect 59878 -5500 59930 -5448
rect 60071 -5500 60123 -5448
rect 60260 -5501 60312 -5449
rect 60454 -5500 60506 -5448
rect 60645 -5500 60697 -5448
rect 60838 -5500 60890 -5448
rect 61030 -5500 61082 -5448
rect 61222 -5501 61274 -5449
rect 61415 -5499 61467 -5447
rect 61605 -5499 61657 -5447
rect 61798 -5501 61850 -5449
rect 61990 -5500 62042 -5448
rect 62183 -5499 62235 -5447
rect 62374 -5499 62426 -5447
rect 62566 -5500 62618 -5448
rect 62757 -5500 62809 -5448
rect 62949 -5500 63001 -5448
rect 63143 -5499 63195 -5447
rect 63335 -5500 63387 -5448
rect 63525 -5501 63577 -5449
rect 63716 -5502 63768 -5450
rect 63909 -5500 63961 -5448
rect 64102 -5499 64154 -5447
rect 64295 -5500 64347 -5448
rect 64486 -5500 64538 -5448
rect 64677 -5500 64729 -5448
rect 64870 -5500 64922 -5448
rect 65063 -5500 65115 -5448
rect 65254 -5500 65306 -5448
rect 65445 -5499 65497 -5447
rect 65636 -5499 65688 -5447
rect 65829 -5500 65881 -5448
rect 66023 -5500 66075 -5448
rect 66211 -5501 66263 -5449
rect 66405 -5509 66457 -5457
rect 49991 -5637 50043 -5585
rect 50182 -5639 50234 -5587
rect 50374 -5638 50426 -5586
rect 50566 -5641 50618 -5589
rect 50760 -5640 50812 -5588
rect 50950 -5640 51002 -5588
rect 51145 -5638 51197 -5586
rect 51336 -5637 51388 -5585
rect 51531 -5639 51583 -5587
rect 51721 -5639 51773 -5587
rect 51911 -5638 51963 -5586
rect 52104 -5637 52156 -5585
rect 52295 -5637 52347 -5585
rect 52491 -5639 52543 -5587
rect 52680 -5639 52732 -5587
rect 52874 -5639 52926 -5587
rect 53063 -5639 53115 -5587
rect 53255 -5640 53307 -5588
rect 53448 -5640 53500 -5588
rect 53639 -5640 53691 -5588
rect 53831 -5639 53883 -5587
rect 54023 -5640 54075 -5588
rect 54216 -5640 54268 -5588
rect 54407 -5640 54459 -5588
rect 54599 -5639 54651 -5587
rect 54792 -5640 54844 -5588
rect 54984 -5640 55036 -5588
rect 55175 -5640 55227 -5588
rect 55366 -5640 55418 -5588
rect 55558 -5640 55610 -5588
rect 55751 -5639 55803 -5587
rect 55942 -5639 55994 -5587
rect 56136 -5640 56188 -5588
rect 56328 -5640 56380 -5588
rect 56520 -5640 56572 -5588
rect 56712 -5640 56764 -5588
rect 56904 -5640 56956 -5588
rect 57096 -5640 57148 -5588
rect 57288 -5640 57340 -5588
rect 57479 -5640 57531 -5588
rect 57671 -5640 57723 -5588
rect 57864 -5640 57916 -5588
rect 58056 -5640 58108 -5588
rect 58248 -5640 58300 -5588
rect 58439 -5640 58491 -5588
rect 58631 -5640 58683 -5588
rect 58822 -5640 58874 -5588
rect 59013 -5640 59065 -5588
rect 59207 -5640 59259 -5588
rect 59399 -5640 59451 -5588
rect 59592 -5639 59644 -5587
rect 59783 -5640 59835 -5588
rect 59975 -5640 60027 -5588
rect 60168 -5640 60220 -5588
rect 60360 -5640 60412 -5588
rect 60553 -5639 60605 -5587
rect 60744 -5640 60796 -5588
rect 60936 -5640 60988 -5588
rect 61127 -5640 61179 -5588
rect 61319 -5640 61371 -5588
rect 61511 -5640 61563 -5588
rect 61704 -5640 61756 -5588
rect 61895 -5640 61947 -5588
rect 62087 -5640 62139 -5588
rect 62279 -5639 62331 -5587
rect 62471 -5640 62523 -5588
rect 62661 -5640 62713 -5588
rect 62855 -5640 62907 -5588
rect 63047 -5639 63099 -5587
rect 63238 -5640 63290 -5588
rect 63431 -5640 63483 -5588
rect 63622 -5639 63674 -5587
rect 63814 -5640 63866 -5588
rect 64005 -5640 64057 -5588
rect 64199 -5639 64251 -5587
rect 64390 -5640 64442 -5588
rect 64582 -5640 64634 -5588
rect 64774 -5640 64826 -5588
rect 64966 -5640 65018 -5588
rect 65159 -5640 65211 -5588
rect 65350 -5640 65402 -5588
rect 65543 -5639 65595 -5587
rect 65734 -5640 65786 -5588
rect 65927 -5640 65979 -5588
rect 66118 -5640 66170 -5588
rect 66309 -5638 66361 -5586
rect 66504 -5640 66556 -5588
rect 49430 -6126 49482 -6074
rect 52047 -6123 52099 -6071
rect 52237 -6122 52289 -6070
rect 52429 -6121 52481 -6069
rect 52620 -6121 52672 -6069
rect 52814 -6121 52866 -6069
rect 53004 -6122 53056 -6070
rect 53198 -6121 53250 -6069
rect 53390 -6121 53442 -6069
rect 53581 -6122 53633 -6070
rect 53776 -6122 53828 -6070
rect 53966 -6122 54018 -6070
rect 54157 -6122 54209 -6070
rect 54349 -6122 54401 -6070
rect 54542 -6121 54594 -6069
rect 54734 -6122 54786 -6070
rect 54926 -6122 54978 -6070
rect 55119 -6122 55171 -6070
rect 55310 -6121 55362 -6069
rect 55502 -6122 55554 -6070
rect 55694 -6121 55746 -6069
rect 55886 -6121 55938 -6069
rect 56077 -6122 56129 -6070
rect 56270 -6121 56322 -6069
rect 56462 -6121 56514 -6069
rect 56656 -6122 56708 -6070
rect 56847 -6123 56899 -6071
rect 57036 -6122 57088 -6070
rect 57229 -6122 57281 -6070
rect 57422 -6122 57474 -6070
rect 57613 -6121 57665 -6069
rect 57804 -6121 57856 -6069
rect 51949 -6262 52001 -6210
rect 52141 -6262 52193 -6210
rect 52334 -6262 52386 -6210
rect 52526 -6262 52578 -6210
rect 52719 -6262 52771 -6210
rect 52911 -6261 52963 -6209
rect 53102 -6262 53154 -6210
rect 53294 -6262 53346 -6210
rect 53486 -6261 53538 -6209
rect 53678 -6261 53730 -6209
rect 53870 -6262 53922 -6210
rect 54062 -6261 54114 -6209
rect 54254 -6262 54306 -6210
rect 54445 -6261 54497 -6209
rect 54639 -6262 54691 -6210
rect 54829 -6262 54881 -6210
rect 55021 -6262 55073 -6210
rect 55214 -6262 55266 -6210
rect 55405 -6262 55457 -6210
rect 55598 -6261 55650 -6209
rect 55791 -6262 55843 -6210
rect 55982 -6262 56034 -6210
rect 56175 -6262 56227 -6210
rect 56365 -6262 56417 -6210
rect 56559 -6261 56611 -6209
rect 56748 -6262 56800 -6210
rect 56941 -6262 56993 -6210
rect 57134 -6262 57186 -6210
rect 57324 -6262 57376 -6210
rect 57517 -6261 57569 -6209
rect 57706 -6261 57758 -6209
rect 51116 -6448 51168 -6396
rect 52040 -6380 52100 -6320
rect 57800 -6370 57860 -6310
rect 66918 -6002 66970 -5950
rect 58241 -6122 58293 -6070
rect 58431 -6121 58483 -6069
rect 58623 -6120 58675 -6068
rect 58814 -6120 58866 -6068
rect 59008 -6120 59060 -6068
rect 59198 -6121 59250 -6069
rect 59392 -6120 59444 -6068
rect 59584 -6120 59636 -6068
rect 59775 -6121 59827 -6069
rect 59970 -6121 60022 -6069
rect 60160 -6121 60212 -6069
rect 60351 -6121 60403 -6069
rect 60543 -6121 60595 -6069
rect 60736 -6120 60788 -6068
rect 60928 -6121 60980 -6069
rect 61120 -6121 61172 -6069
rect 61313 -6121 61365 -6069
rect 61504 -6120 61556 -6068
rect 61696 -6121 61748 -6069
rect 61888 -6120 61940 -6068
rect 62080 -6120 62132 -6068
rect 62271 -6121 62323 -6069
rect 62464 -6120 62516 -6068
rect 62656 -6120 62708 -6068
rect 62850 -6121 62902 -6069
rect 63041 -6122 63093 -6070
rect 63230 -6121 63282 -6069
rect 63423 -6121 63475 -6069
rect 63616 -6121 63668 -6069
rect 63807 -6120 63859 -6068
rect 63998 -6120 64050 -6068
rect 58143 -6261 58195 -6209
rect 58335 -6261 58387 -6209
rect 58528 -6261 58580 -6209
rect 58720 -6261 58772 -6209
rect 58913 -6261 58965 -6209
rect 59105 -6260 59157 -6208
rect 59296 -6261 59348 -6209
rect 59488 -6261 59540 -6209
rect 59680 -6260 59732 -6208
rect 59872 -6260 59924 -6208
rect 60064 -6261 60116 -6209
rect 60256 -6260 60308 -6208
rect 60448 -6261 60500 -6209
rect 60639 -6260 60691 -6208
rect 60833 -6261 60885 -6209
rect 61023 -6261 61075 -6209
rect 61215 -6261 61267 -6209
rect 61408 -6261 61460 -6209
rect 61599 -6261 61651 -6209
rect 61792 -6260 61844 -6208
rect 61985 -6261 62037 -6209
rect 62176 -6261 62228 -6209
rect 62369 -6261 62421 -6209
rect 62559 -6261 62611 -6209
rect 62753 -6260 62805 -6208
rect 62942 -6261 62994 -6209
rect 63135 -6261 63187 -6209
rect 63328 -6261 63380 -6209
rect 63518 -6261 63570 -6209
rect 63711 -6260 63763 -6208
rect 63900 -6260 63952 -6208
rect 68930 -6272 69296 -5188
rect 58230 -6370 58290 -6310
rect 63990 -6360 64050 -6300
rect 64530 -6432 64582 -6380
rect 51116 -6552 51168 -6500
rect 64536 -6548 64588 -6496
rect 47254 -7752 47614 -6678
rect 49436 -6924 49488 -6872
rect 52048 -6741 52100 -6689
rect 52238 -6740 52290 -6688
rect 52430 -6739 52482 -6687
rect 52621 -6739 52673 -6687
rect 52815 -6739 52867 -6687
rect 53005 -6740 53057 -6688
rect 53199 -6739 53251 -6687
rect 53391 -6739 53443 -6687
rect 53582 -6740 53634 -6688
rect 53777 -6740 53829 -6688
rect 53967 -6740 54019 -6688
rect 54158 -6740 54210 -6688
rect 54350 -6740 54402 -6688
rect 54543 -6739 54595 -6687
rect 54735 -6740 54787 -6688
rect 54927 -6740 54979 -6688
rect 55120 -6740 55172 -6688
rect 55311 -6739 55363 -6687
rect 55503 -6740 55555 -6688
rect 55695 -6739 55747 -6687
rect 55887 -6739 55939 -6687
rect 56078 -6740 56130 -6688
rect 56271 -6739 56323 -6687
rect 56463 -6739 56515 -6687
rect 56657 -6740 56709 -6688
rect 56848 -6741 56900 -6689
rect 57037 -6740 57089 -6688
rect 57230 -6740 57282 -6688
rect 57423 -6740 57475 -6688
rect 57614 -6739 57666 -6687
rect 57805 -6739 57857 -6687
rect 51950 -6880 52002 -6828
rect 52142 -6880 52194 -6828
rect 52335 -6880 52387 -6828
rect 52527 -6880 52579 -6828
rect 52720 -6880 52772 -6828
rect 52912 -6879 52964 -6827
rect 53103 -6880 53155 -6828
rect 53295 -6880 53347 -6828
rect 53487 -6879 53539 -6827
rect 53679 -6879 53731 -6827
rect 53871 -6880 53923 -6828
rect 54063 -6879 54115 -6827
rect 54255 -6880 54307 -6828
rect 54446 -6879 54498 -6827
rect 54640 -6880 54692 -6828
rect 54830 -6880 54882 -6828
rect 55022 -6880 55074 -6828
rect 55215 -6880 55267 -6828
rect 55406 -6880 55458 -6828
rect 55599 -6879 55651 -6827
rect 55792 -6880 55844 -6828
rect 55983 -6880 56035 -6828
rect 56176 -6880 56228 -6828
rect 56366 -6880 56418 -6828
rect 56560 -6879 56612 -6827
rect 56749 -6880 56801 -6828
rect 56942 -6880 56994 -6828
rect 57135 -6880 57187 -6828
rect 57325 -6880 57377 -6828
rect 57518 -6879 57570 -6827
rect 57707 -6879 57759 -6827
rect 58236 -6740 58288 -6688
rect 58426 -6739 58478 -6687
rect 58618 -6738 58670 -6686
rect 58809 -6738 58861 -6686
rect 59003 -6738 59055 -6686
rect 59193 -6739 59245 -6687
rect 59387 -6738 59439 -6686
rect 59579 -6738 59631 -6686
rect 59770 -6739 59822 -6687
rect 59965 -6739 60017 -6687
rect 60155 -6739 60207 -6687
rect 60346 -6739 60398 -6687
rect 60538 -6739 60590 -6687
rect 60731 -6738 60783 -6686
rect 60923 -6739 60975 -6687
rect 61115 -6739 61167 -6687
rect 61308 -6739 61360 -6687
rect 61499 -6738 61551 -6686
rect 61691 -6739 61743 -6687
rect 61883 -6738 61935 -6686
rect 62075 -6738 62127 -6686
rect 62266 -6739 62318 -6687
rect 62459 -6738 62511 -6686
rect 62651 -6738 62703 -6686
rect 62845 -6739 62897 -6687
rect 63036 -6740 63088 -6688
rect 63225 -6739 63277 -6687
rect 63418 -6739 63470 -6687
rect 63611 -6739 63663 -6687
rect 63802 -6738 63854 -6686
rect 63993 -6738 64045 -6686
rect 58138 -6879 58190 -6827
rect 58330 -6879 58382 -6827
rect 58523 -6879 58575 -6827
rect 58715 -6879 58767 -6827
rect 58908 -6879 58960 -6827
rect 59100 -6878 59152 -6826
rect 59291 -6879 59343 -6827
rect 59483 -6879 59535 -6827
rect 59675 -6878 59727 -6826
rect 59867 -6878 59919 -6826
rect 60059 -6879 60111 -6827
rect 60251 -6878 60303 -6826
rect 60443 -6879 60495 -6827
rect 60634 -6878 60686 -6826
rect 60828 -6879 60880 -6827
rect 61018 -6879 61070 -6827
rect 61210 -6879 61262 -6827
rect 61403 -6879 61455 -6827
rect 61594 -6879 61646 -6827
rect 61787 -6878 61839 -6826
rect 61980 -6879 62032 -6827
rect 62171 -6879 62223 -6827
rect 62364 -6879 62416 -6827
rect 62554 -6879 62606 -6827
rect 62748 -6878 62800 -6826
rect 62937 -6879 62989 -6827
rect 63130 -6879 63182 -6827
rect 63323 -6879 63375 -6827
rect 63513 -6879 63565 -6827
rect 63706 -6878 63758 -6826
rect 63895 -6878 63947 -6826
rect 66912 -6902 66964 -6850
rect 50087 -7354 50139 -7302
rect 50277 -7353 50329 -7301
rect 50470 -7356 50522 -7304
rect 50662 -7351 50714 -7299
rect 50854 -7355 50906 -7303
rect 51046 -7350 51098 -7298
rect 51238 -7351 51290 -7299
rect 51428 -7350 51480 -7298
rect 51622 -7361 51674 -7309
rect 51811 -7359 51863 -7307
rect 52001 -7359 52053 -7307
rect 52200 -7360 52252 -7308
rect 52392 -7359 52444 -7307
rect 52582 -7360 52634 -7308
rect 52774 -7353 52826 -7301
rect 52966 -7355 53018 -7303
rect 53159 -7354 53211 -7302
rect 53351 -7352 53403 -7300
rect 53542 -7352 53594 -7300
rect 53736 -7357 53788 -7305
rect 53927 -7353 53979 -7301
rect 54119 -7349 54171 -7297
rect 54312 -7353 54364 -7301
rect 54504 -7353 54556 -7301
rect 54697 -7354 54749 -7302
rect 54889 -7352 54941 -7300
rect 55080 -7351 55132 -7299
rect 55271 -7350 55323 -7298
rect 55464 -7350 55516 -7298
rect 55655 -7359 55707 -7307
rect 55846 -7360 55898 -7308
rect 56036 -7361 56088 -7309
rect 56230 -7365 56282 -7313
rect 56422 -7367 56474 -7315
rect 56616 -7366 56668 -7314
rect 56808 -7363 56860 -7311
rect 56997 -7360 57049 -7308
rect 57191 -7358 57243 -7306
rect 57384 -7359 57436 -7307
rect 57577 -7360 57629 -7308
rect 57766 -7360 57818 -7308
rect 57959 -7360 58011 -7308
rect 58151 -7360 58203 -7308
rect 58342 -7360 58394 -7308
rect 58535 -7360 58587 -7308
rect 58726 -7359 58778 -7307
rect 58921 -7360 58973 -7308
rect 59110 -7360 59162 -7308
rect 59303 -7360 59355 -7308
rect 59495 -7360 59547 -7308
rect 59686 -7360 59738 -7308
rect 59878 -7360 59930 -7308
rect 60071 -7360 60123 -7308
rect 60260 -7361 60312 -7309
rect 60454 -7360 60506 -7308
rect 60645 -7360 60697 -7308
rect 60838 -7360 60890 -7308
rect 61030 -7360 61082 -7308
rect 61222 -7361 61274 -7309
rect 61415 -7359 61467 -7307
rect 61605 -7359 61657 -7307
rect 61798 -7361 61850 -7309
rect 61990 -7360 62042 -7308
rect 62183 -7359 62235 -7307
rect 62374 -7359 62426 -7307
rect 62566 -7360 62618 -7308
rect 62757 -7360 62809 -7308
rect 62949 -7360 63001 -7308
rect 63143 -7359 63195 -7307
rect 63335 -7360 63387 -7308
rect 63525 -7361 63577 -7309
rect 63716 -7362 63768 -7310
rect 63909 -7360 63961 -7308
rect 64102 -7359 64154 -7307
rect 64295 -7360 64347 -7308
rect 64486 -7360 64538 -7308
rect 64677 -7360 64729 -7308
rect 64870 -7360 64922 -7308
rect 65063 -7360 65115 -7308
rect 65254 -7360 65306 -7308
rect 65445 -7359 65497 -7307
rect 65636 -7359 65688 -7307
rect 65829 -7360 65881 -7308
rect 66023 -7360 66075 -7308
rect 66211 -7361 66263 -7309
rect 66405 -7369 66457 -7317
rect 49991 -7497 50043 -7445
rect 50182 -7499 50234 -7447
rect 50374 -7498 50426 -7446
rect 50566 -7501 50618 -7449
rect 50760 -7500 50812 -7448
rect 50950 -7500 51002 -7448
rect 51145 -7498 51197 -7446
rect 51336 -7497 51388 -7445
rect 51531 -7499 51583 -7447
rect 51721 -7499 51773 -7447
rect 51911 -7498 51963 -7446
rect 52104 -7497 52156 -7445
rect 52295 -7497 52347 -7445
rect 52491 -7499 52543 -7447
rect 52680 -7499 52732 -7447
rect 52874 -7499 52926 -7447
rect 53063 -7499 53115 -7447
rect 53255 -7500 53307 -7448
rect 53448 -7500 53500 -7448
rect 53639 -7500 53691 -7448
rect 53831 -7499 53883 -7447
rect 54023 -7500 54075 -7448
rect 54216 -7500 54268 -7448
rect 54407 -7500 54459 -7448
rect 54599 -7499 54651 -7447
rect 54792 -7500 54844 -7448
rect 54984 -7500 55036 -7448
rect 55175 -7500 55227 -7448
rect 55366 -7500 55418 -7448
rect 55558 -7500 55610 -7448
rect 55751 -7499 55803 -7447
rect 55942 -7499 55994 -7447
rect 56136 -7500 56188 -7448
rect 56328 -7500 56380 -7448
rect 56520 -7500 56572 -7448
rect 56712 -7500 56764 -7448
rect 56904 -7500 56956 -7448
rect 57096 -7500 57148 -7448
rect 57288 -7500 57340 -7448
rect 57479 -7500 57531 -7448
rect 57671 -7500 57723 -7448
rect 57864 -7500 57916 -7448
rect 58056 -7500 58108 -7448
rect 58248 -7500 58300 -7448
rect 58439 -7500 58491 -7448
rect 58631 -7500 58683 -7448
rect 58822 -7500 58874 -7448
rect 59013 -7500 59065 -7448
rect 59207 -7500 59259 -7448
rect 59399 -7500 59451 -7448
rect 59592 -7499 59644 -7447
rect 59783 -7500 59835 -7448
rect 59975 -7500 60027 -7448
rect 60168 -7500 60220 -7448
rect 60360 -7500 60412 -7448
rect 60553 -7499 60605 -7447
rect 60744 -7500 60796 -7448
rect 60936 -7500 60988 -7448
rect 61127 -7500 61179 -7448
rect 61319 -7500 61371 -7448
rect 61511 -7500 61563 -7448
rect 61704 -7500 61756 -7448
rect 61895 -7500 61947 -7448
rect 62087 -7500 62139 -7448
rect 62279 -7499 62331 -7447
rect 62471 -7500 62523 -7448
rect 62661 -7500 62713 -7448
rect 62855 -7500 62907 -7448
rect 63047 -7499 63099 -7447
rect 63238 -7500 63290 -7448
rect 63431 -7500 63483 -7448
rect 63622 -7499 63674 -7447
rect 63814 -7500 63866 -7448
rect 64005 -7500 64057 -7448
rect 64199 -7499 64251 -7447
rect 64390 -7500 64442 -7448
rect 64582 -7500 64634 -7448
rect 64774 -7500 64826 -7448
rect 64966 -7500 65018 -7448
rect 65159 -7500 65211 -7448
rect 65350 -7500 65402 -7448
rect 65543 -7499 65595 -7447
rect 65734 -7500 65786 -7448
rect 65927 -7500 65979 -7448
rect 66118 -7500 66170 -7448
rect 66309 -7498 66361 -7446
rect 66504 -7500 66556 -7448
rect 48274 -7764 48446 -7706
rect 49940 -7756 66588 -7664
rect 68120 -7768 68292 -7710
rect 68924 -7756 69290 -6672
<< metal2 >>
rect 68894 -4738 69326 -4736
rect 68674 -4740 69326 -4738
rect 47224 -5130 69326 -4740
rect 47224 -5190 47652 -5130
rect 47224 -6264 47260 -5190
rect 47620 -6264 47652 -5190
rect 48286 -5178 48458 -5168
rect 68070 -5178 68242 -5168
rect 48286 -5246 48458 -5236
rect 49920 -5188 66568 -5178
rect 68070 -5246 68242 -5236
rect 68894 -5188 69326 -5130
rect 49920 -5290 66568 -5280
rect 50090 -5432 50160 -5290
rect 50087 -5440 50160 -5432
rect 50277 -5440 50329 -5431
rect 50470 -5440 50522 -5434
rect 50662 -5439 50714 -5430
rect 50087 -5441 50662 -5440
rect 50087 -5442 50277 -5441
rect 50139 -5470 50277 -5442
rect 50087 -5504 50139 -5494
rect 50329 -5444 50662 -5441
rect 50329 -5470 50470 -5444
rect 50277 -5503 50329 -5493
rect 50522 -5470 50662 -5444
rect 50470 -5506 50522 -5496
rect 50854 -5440 50906 -5433
rect 51046 -5438 51098 -5430
rect 50714 -5443 51046 -5440
rect 50714 -5470 50854 -5443
rect 50662 -5501 50714 -5491
rect 50906 -5470 51046 -5443
rect 50854 -5505 50906 -5495
rect 51238 -5439 51290 -5430
rect 51098 -5470 51238 -5440
rect 51046 -5500 51098 -5490
rect 51428 -5438 51480 -5430
rect 51290 -5470 51428 -5440
rect 51238 -5501 51290 -5491
rect 51622 -5440 51674 -5439
rect 51811 -5440 51863 -5437
rect 52001 -5440 52053 -5437
rect 52200 -5440 52252 -5438
rect 52392 -5440 52444 -5437
rect 52582 -5440 52634 -5438
rect 52774 -5440 52826 -5431
rect 52966 -5440 53018 -5433
rect 53159 -5440 53211 -5432
rect 53351 -5440 53403 -5430
rect 53542 -5440 53594 -5430
rect 53736 -5440 53788 -5435
rect 53927 -5440 53979 -5431
rect 54119 -5437 54171 -5430
rect 51480 -5441 53351 -5440
rect 51480 -5447 52774 -5441
rect 51480 -5449 51811 -5447
rect 51480 -5470 51622 -5449
rect 51428 -5500 51480 -5490
rect 51674 -5470 51811 -5449
rect 51622 -5511 51674 -5501
rect 51863 -5470 52001 -5447
rect 51811 -5509 51863 -5499
rect 52053 -5448 52392 -5447
rect 52053 -5470 52200 -5448
rect 52001 -5509 52053 -5499
rect 52252 -5470 52392 -5448
rect 52200 -5510 52252 -5500
rect 52444 -5448 52774 -5447
rect 52444 -5470 52582 -5448
rect 52392 -5509 52444 -5499
rect 52634 -5470 52774 -5448
rect 52582 -5510 52634 -5500
rect 52826 -5442 53351 -5441
rect 52826 -5443 53159 -5442
rect 52826 -5470 52966 -5443
rect 52774 -5503 52826 -5493
rect 53018 -5470 53159 -5443
rect 52966 -5505 53018 -5495
rect 53211 -5470 53351 -5442
rect 53159 -5504 53211 -5494
rect 53403 -5470 53542 -5440
rect 53351 -5502 53403 -5492
rect 53594 -5441 54119 -5440
rect 53594 -5445 53927 -5441
rect 53594 -5470 53736 -5445
rect 53542 -5502 53594 -5492
rect 53788 -5470 53927 -5445
rect 53736 -5507 53788 -5497
rect 53979 -5470 54119 -5441
rect 53927 -5503 53979 -5493
rect 54312 -5440 54364 -5431
rect 54504 -5440 54556 -5431
rect 54697 -5440 54749 -5432
rect 54889 -5440 54941 -5430
rect 55080 -5439 55132 -5430
rect 54171 -5441 54889 -5440
rect 54171 -5470 54312 -5441
rect 54119 -5499 54171 -5489
rect 54364 -5470 54504 -5441
rect 54312 -5503 54364 -5493
rect 54556 -5442 54889 -5441
rect 54556 -5470 54697 -5442
rect 54504 -5503 54556 -5493
rect 54749 -5470 54889 -5442
rect 54697 -5504 54749 -5494
rect 54941 -5470 55080 -5440
rect 54889 -5502 54941 -5492
rect 55271 -5438 55323 -5430
rect 55132 -5470 55271 -5440
rect 55080 -5501 55132 -5491
rect 55464 -5438 55516 -5430
rect 55323 -5470 55464 -5440
rect 55271 -5500 55323 -5490
rect 55655 -5440 55707 -5437
rect 55846 -5440 55898 -5438
rect 56036 -5440 56088 -5439
rect 56997 -5440 57049 -5438
rect 57191 -5440 57243 -5436
rect 57384 -5440 57436 -5437
rect 57577 -5440 57629 -5438
rect 57766 -5440 57818 -5438
rect 57959 -5440 58011 -5438
rect 58151 -5440 58203 -5438
rect 58342 -5440 58394 -5438
rect 58535 -5440 58587 -5438
rect 58726 -5440 58778 -5437
rect 58921 -5440 58973 -5438
rect 59110 -5440 59162 -5438
rect 59303 -5440 59355 -5438
rect 59495 -5440 59547 -5438
rect 59686 -5440 59738 -5438
rect 59878 -5440 59930 -5438
rect 60071 -5440 60123 -5438
rect 60260 -5440 60312 -5439
rect 60454 -5440 60506 -5438
rect 60645 -5440 60697 -5438
rect 60838 -5440 60890 -5438
rect 61030 -5440 61082 -5438
rect 61222 -5440 61274 -5439
rect 61415 -5440 61467 -5437
rect 61605 -5440 61657 -5437
rect 61798 -5440 61850 -5439
rect 61990 -5440 62042 -5438
rect 62183 -5440 62235 -5437
rect 62374 -5440 62426 -5437
rect 62566 -5440 62618 -5438
rect 62757 -5440 62809 -5438
rect 62949 -5440 63001 -5438
rect 63143 -5440 63195 -5437
rect 63335 -5440 63387 -5438
rect 63525 -5440 63577 -5439
rect 63909 -5440 63961 -5438
rect 64102 -5440 64154 -5437
rect 64295 -5440 64347 -5438
rect 64486 -5440 64538 -5438
rect 64677 -5440 64729 -5438
rect 64870 -5440 64922 -5438
rect 65063 -5440 65115 -5438
rect 65254 -5440 65306 -5438
rect 65445 -5440 65497 -5437
rect 65636 -5440 65688 -5437
rect 65829 -5440 65881 -5438
rect 66023 -5440 66075 -5438
rect 66211 -5440 66263 -5439
rect 66400 -5440 66470 -5290
rect 55516 -5446 66470 -5440
rect 55516 -5447 57191 -5446
rect 55516 -5470 55655 -5447
rect 55464 -5500 55516 -5490
rect 55707 -5448 57191 -5447
rect 55707 -5470 55846 -5448
rect 55655 -5509 55707 -5499
rect 55898 -5449 56997 -5448
rect 55898 -5470 56036 -5449
rect 55846 -5510 55898 -5500
rect 56088 -5451 56997 -5449
rect 56088 -5453 56808 -5451
rect 56088 -5470 56230 -5453
rect 56036 -5511 56088 -5501
rect 56282 -5454 56808 -5453
rect 56282 -5455 56616 -5454
rect 56282 -5470 56422 -5455
rect 56230 -5515 56282 -5505
rect 56474 -5470 56616 -5455
rect 56422 -5517 56474 -5507
rect 56668 -5470 56808 -5454
rect 56616 -5516 56668 -5506
rect 56860 -5470 56997 -5451
rect 56808 -5513 56860 -5503
rect 57049 -5470 57191 -5448
rect 56997 -5510 57049 -5500
rect 57243 -5447 66470 -5446
rect 57243 -5470 57384 -5447
rect 57191 -5508 57243 -5498
rect 57436 -5448 58726 -5447
rect 57436 -5470 57577 -5448
rect 57384 -5509 57436 -5499
rect 57629 -5470 57766 -5448
rect 57577 -5510 57629 -5500
rect 57818 -5470 57959 -5448
rect 57766 -5510 57818 -5500
rect 58011 -5470 58151 -5448
rect 57959 -5510 58011 -5500
rect 58203 -5470 58342 -5448
rect 58151 -5510 58203 -5500
rect 58394 -5470 58535 -5448
rect 58342 -5510 58394 -5500
rect 58587 -5470 58726 -5448
rect 58535 -5510 58587 -5500
rect 58778 -5448 61415 -5447
rect 58778 -5470 58921 -5448
rect 58726 -5509 58778 -5499
rect 58973 -5470 59110 -5448
rect 58921 -5510 58973 -5500
rect 59162 -5470 59303 -5448
rect 59110 -5510 59162 -5500
rect 59355 -5470 59495 -5448
rect 59303 -5510 59355 -5500
rect 59547 -5470 59686 -5448
rect 59495 -5510 59547 -5500
rect 59738 -5470 59878 -5448
rect 59686 -5510 59738 -5500
rect 59930 -5470 60071 -5448
rect 59878 -5510 59930 -5500
rect 60123 -5449 60454 -5448
rect 60123 -5470 60260 -5449
rect 60071 -5510 60123 -5500
rect 60312 -5470 60454 -5449
rect 60260 -5511 60312 -5501
rect 60506 -5470 60645 -5448
rect 60454 -5510 60506 -5500
rect 60697 -5470 60838 -5448
rect 60645 -5510 60697 -5500
rect 60890 -5470 61030 -5448
rect 60838 -5510 60890 -5500
rect 61082 -5449 61415 -5448
rect 61082 -5470 61222 -5449
rect 61030 -5510 61082 -5500
rect 61274 -5470 61415 -5449
rect 61222 -5511 61274 -5501
rect 61467 -5470 61605 -5447
rect 61415 -5509 61467 -5499
rect 61657 -5448 62183 -5447
rect 61657 -5449 61990 -5448
rect 61657 -5470 61798 -5449
rect 61605 -5509 61657 -5499
rect 61850 -5470 61990 -5449
rect 61798 -5511 61850 -5501
rect 62042 -5470 62183 -5448
rect 61990 -5510 62042 -5500
rect 62235 -5470 62374 -5447
rect 62183 -5509 62235 -5499
rect 62426 -5448 63143 -5447
rect 62426 -5470 62566 -5448
rect 62374 -5509 62426 -5499
rect 62618 -5470 62757 -5448
rect 62566 -5510 62618 -5500
rect 62809 -5470 62949 -5448
rect 62757 -5510 62809 -5500
rect 63001 -5470 63143 -5448
rect 62949 -5510 63001 -5500
rect 63195 -5448 64102 -5447
rect 63195 -5470 63335 -5448
rect 63143 -5509 63195 -5499
rect 63387 -5449 63909 -5448
rect 63387 -5470 63525 -5449
rect 63335 -5510 63387 -5500
rect 63577 -5450 63909 -5449
rect 63577 -5470 63716 -5450
rect 63525 -5511 63577 -5501
rect 63768 -5470 63909 -5450
rect 63716 -5512 63768 -5502
rect 63961 -5470 64102 -5448
rect 63909 -5510 63961 -5500
rect 64154 -5448 65445 -5447
rect 64154 -5470 64295 -5448
rect 64102 -5509 64154 -5499
rect 64347 -5470 64486 -5448
rect 64295 -5510 64347 -5500
rect 64538 -5470 64677 -5448
rect 64486 -5510 64538 -5500
rect 64729 -5470 64870 -5448
rect 64677 -5510 64729 -5500
rect 64922 -5470 65063 -5448
rect 64870 -5510 64922 -5500
rect 65115 -5470 65254 -5448
rect 65063 -5510 65115 -5500
rect 65306 -5470 65445 -5448
rect 65254 -5510 65306 -5500
rect 65497 -5470 65636 -5447
rect 65445 -5509 65497 -5499
rect 65688 -5448 66470 -5447
rect 65688 -5470 65829 -5448
rect 65636 -5509 65688 -5499
rect 65881 -5470 66023 -5448
rect 65829 -5510 65881 -5500
rect 66075 -5449 66470 -5448
rect 66075 -5470 66211 -5449
rect 66023 -5510 66075 -5500
rect 66263 -5457 66470 -5449
rect 66263 -5470 66405 -5457
rect 66211 -5511 66263 -5501
rect 66457 -5470 66470 -5457
rect 66405 -5519 66457 -5509
rect 49991 -5585 50043 -5575
rect 50182 -5587 50234 -5577
rect 50043 -5630 50182 -5600
rect 49991 -5647 50043 -5637
rect 50374 -5586 50426 -5576
rect 50234 -5630 50374 -5600
rect 50182 -5649 50234 -5639
rect 50566 -5589 50618 -5579
rect 50426 -5630 50566 -5600
rect 50374 -5648 50426 -5638
rect 50760 -5588 50812 -5578
rect 50618 -5630 50760 -5600
rect 50566 -5651 50618 -5641
rect 50950 -5588 51002 -5578
rect 50812 -5630 50950 -5600
rect 50760 -5650 50812 -5640
rect 51145 -5586 51197 -5576
rect 51002 -5630 51145 -5600
rect 50950 -5650 51002 -5640
rect 51336 -5585 51388 -5575
rect 51197 -5630 51336 -5600
rect 51145 -5648 51197 -5638
rect 51531 -5587 51583 -5577
rect 51388 -5630 51531 -5600
rect 51336 -5647 51388 -5637
rect 51721 -5587 51773 -5577
rect 51583 -5630 51721 -5600
rect 51531 -5649 51583 -5639
rect 51911 -5586 51963 -5576
rect 51773 -5630 51911 -5600
rect 51721 -5649 51773 -5639
rect 52104 -5585 52156 -5575
rect 51963 -5630 52104 -5600
rect 51911 -5648 51963 -5638
rect 52050 -5637 52104 -5630
rect 52295 -5585 52347 -5575
rect 52156 -5630 52295 -5600
rect 52050 -5647 52156 -5637
rect 52491 -5587 52543 -5577
rect 52347 -5630 52491 -5600
rect 52295 -5647 52347 -5637
rect 52430 -5639 52491 -5630
rect 52680 -5587 52732 -5577
rect 52543 -5630 52680 -5600
rect 52050 -6060 52110 -5647
rect 52430 -5649 52543 -5639
rect 52874 -5587 52926 -5577
rect 52732 -5630 52874 -5600
rect 52680 -5649 52732 -5639
rect 52820 -5639 52874 -5630
rect 53063 -5587 53115 -5577
rect 52926 -5630 53063 -5600
rect 52820 -5649 52926 -5639
rect 53255 -5588 53307 -5578
rect 53115 -5630 53255 -5600
rect 53063 -5649 53115 -5639
rect 53200 -5640 53255 -5630
rect 53448 -5588 53500 -5578
rect 53307 -5630 53448 -5600
rect 52430 -6059 52490 -5649
rect 52820 -6059 52880 -5649
rect 53200 -5650 53307 -5640
rect 53639 -5588 53691 -5578
rect 53500 -5630 53639 -5600
rect 53448 -5650 53500 -5640
rect 53580 -5640 53639 -5630
rect 53831 -5587 53883 -5577
rect 53691 -5630 53831 -5600
rect 53580 -5650 53691 -5640
rect 54023 -5588 54075 -5578
rect 53883 -5630 54023 -5600
rect 53831 -5649 53883 -5639
rect 53970 -5640 54023 -5630
rect 54216 -5588 54268 -5578
rect 54075 -5630 54216 -5600
rect 53970 -5650 54075 -5640
rect 54407 -5588 54459 -5578
rect 54268 -5630 54407 -5600
rect 54216 -5650 54268 -5640
rect 54350 -5640 54407 -5630
rect 54599 -5587 54651 -5577
rect 54459 -5630 54599 -5600
rect 54350 -5650 54459 -5640
rect 54792 -5588 54844 -5578
rect 54651 -5630 54792 -5600
rect 54599 -5649 54651 -5639
rect 54740 -5640 54792 -5630
rect 54984 -5588 55036 -5578
rect 54844 -5630 54984 -5600
rect 54740 -5650 54844 -5640
rect 55175 -5588 55227 -5578
rect 55036 -5630 55175 -5600
rect 54984 -5650 55036 -5640
rect 55120 -5640 55175 -5630
rect 55366 -5588 55418 -5578
rect 55227 -5630 55366 -5600
rect 55120 -5650 55227 -5640
rect 55558 -5588 55610 -5578
rect 55418 -5630 55558 -5600
rect 55366 -5650 55418 -5640
rect 55500 -5640 55558 -5630
rect 55751 -5587 55803 -5577
rect 55610 -5630 55751 -5600
rect 55500 -5650 55610 -5640
rect 55942 -5587 55994 -5577
rect 55803 -5630 55942 -5600
rect 55751 -5649 55803 -5639
rect 55890 -5639 55942 -5630
rect 56136 -5588 56188 -5578
rect 55994 -5630 56136 -5600
rect 55890 -5649 55994 -5639
rect 56328 -5588 56380 -5578
rect 56188 -5630 56328 -5600
rect 53200 -6059 53260 -5650
rect 52429 -6060 52490 -6059
rect 52620 -6060 52672 -6059
rect 52814 -6060 52880 -6059
rect 53198 -6060 53260 -6059
rect 53390 -6060 53442 -6059
rect 53580 -6060 53640 -5650
rect 53970 -6060 54030 -5650
rect 54350 -6060 54410 -5650
rect 54542 -6060 54594 -6059
rect 54740 -6060 54800 -5650
rect 55120 -6060 55180 -5650
rect 55310 -6060 55362 -6059
rect 55500 -6060 55560 -5650
rect 55890 -6059 55950 -5649
rect 56136 -5650 56188 -5640
rect 56270 -5640 56328 -5630
rect 56520 -5588 56572 -5578
rect 56380 -5630 56520 -5600
rect 56270 -5650 56380 -5640
rect 56712 -5588 56764 -5578
rect 56572 -5630 56712 -5600
rect 56520 -5650 56572 -5640
rect 56660 -5640 56712 -5630
rect 56904 -5588 56956 -5578
rect 56764 -5630 56904 -5600
rect 56660 -5650 56764 -5640
rect 57096 -5588 57148 -5578
rect 56956 -5630 57096 -5600
rect 56904 -5650 56956 -5640
rect 57040 -5640 57096 -5630
rect 57288 -5588 57340 -5578
rect 57148 -5630 57288 -5600
rect 57040 -5650 57148 -5640
rect 57479 -5588 57531 -5578
rect 57340 -5630 57479 -5600
rect 57288 -5650 57340 -5640
rect 57420 -5640 57479 -5630
rect 57671 -5588 57723 -5578
rect 57531 -5630 57671 -5600
rect 57420 -5650 57531 -5640
rect 57864 -5588 57916 -5578
rect 57723 -5630 57864 -5600
rect 57671 -5650 57723 -5640
rect 57810 -5640 57864 -5630
rect 58056 -5588 58108 -5578
rect 57916 -5630 58056 -5600
rect 57810 -5650 57916 -5640
rect 58248 -5588 58300 -5578
rect 58108 -5630 58248 -5600
rect 58056 -5650 58108 -5640
rect 58240 -5640 58248 -5630
rect 58439 -5588 58491 -5578
rect 58300 -5630 58439 -5600
rect 55694 -6060 55746 -6059
rect 55886 -6060 55950 -6059
rect 56270 -6060 56330 -5650
rect 56462 -6060 56514 -6059
rect 56660 -6060 56720 -5650
rect 57040 -6060 57100 -5650
rect 57420 -6060 57480 -5650
rect 57810 -6059 57870 -5650
rect 57613 -6060 57665 -6059
rect 57804 -6060 57870 -6059
rect 58240 -6060 58300 -5640
rect 58631 -5588 58683 -5578
rect 58491 -5630 58631 -5600
rect 58439 -5650 58491 -5640
rect 58620 -5640 58631 -5630
rect 58822 -5588 58874 -5578
rect 58683 -5630 58822 -5600
rect 58620 -5650 58683 -5640
rect 59013 -5588 59065 -5578
rect 58874 -5630 59013 -5600
rect 58822 -5650 58874 -5640
rect 59010 -5640 59013 -5630
rect 59207 -5588 59259 -5578
rect 59065 -5630 59207 -5600
rect 59065 -5640 59070 -5630
rect 52050 -6061 58300 -6060
rect 58431 -6061 58483 -6059
rect 58620 -6061 58680 -5650
rect 59010 -6058 59070 -5640
rect 59399 -5588 59451 -5578
rect 59259 -5630 59399 -5600
rect 59207 -5650 59259 -5640
rect 59592 -5587 59644 -5577
rect 59451 -5630 59592 -5600
rect 59451 -5640 59460 -5630
rect 59399 -5650 59460 -5640
rect 59783 -5588 59835 -5578
rect 59644 -5630 59783 -5600
rect 59592 -5649 59644 -5639
rect 59780 -5640 59783 -5630
rect 59975 -5588 60027 -5578
rect 59835 -5630 59975 -5600
rect 59835 -5640 59840 -5630
rect 59400 -6058 59460 -5650
rect 58814 -6061 58866 -6058
rect 59008 -6061 59070 -6058
rect 59198 -6061 59250 -6059
rect 59392 -6061 59460 -6058
rect 59584 -6061 59636 -6058
rect 59780 -6059 59840 -5640
rect 60168 -5588 60220 -5578
rect 60027 -5630 60168 -5600
rect 59975 -5650 60027 -5640
rect 60160 -5640 60168 -5630
rect 60360 -5588 60412 -5578
rect 60220 -5630 60360 -5600
rect 59775 -6061 59840 -6059
rect 59970 -6061 60022 -6059
rect 60160 -6061 60220 -5640
rect 60553 -5587 60605 -5577
rect 60412 -5630 60553 -5600
rect 60360 -5650 60412 -5640
rect 60540 -5639 60553 -5630
rect 60744 -5588 60796 -5578
rect 60605 -5630 60744 -5600
rect 60540 -5649 60605 -5639
rect 60936 -5588 60988 -5578
rect 60796 -5630 60936 -5600
rect 60351 -6061 60403 -6059
rect 60540 -6061 60600 -5649
rect 60744 -5650 60796 -5640
rect 60930 -5640 60936 -5630
rect 61127 -5588 61179 -5578
rect 60988 -5630 61127 -5600
rect 60988 -5640 60990 -5630
rect 60736 -6061 60788 -6058
rect 60930 -6059 60990 -5640
rect 61319 -5588 61371 -5578
rect 61179 -5630 61319 -5600
rect 61127 -5650 61179 -5640
rect 61511 -5588 61563 -5578
rect 61371 -5630 61511 -5600
rect 61371 -5640 61380 -5630
rect 61319 -5650 61380 -5640
rect 61704 -5588 61756 -5578
rect 61563 -5630 61704 -5600
rect 61511 -5650 61563 -5640
rect 61700 -5640 61704 -5630
rect 61895 -5588 61947 -5578
rect 61756 -5630 61895 -5600
rect 61756 -5640 61760 -5630
rect 61320 -6059 61380 -5650
rect 60928 -6061 60990 -6059
rect 61120 -6061 61172 -6059
rect 61313 -6061 61380 -6059
rect 61504 -6061 61556 -6058
rect 61700 -6059 61760 -5640
rect 62087 -5588 62139 -5578
rect 61947 -5630 62087 -5600
rect 61895 -5650 61947 -5640
rect 62080 -5640 62087 -5630
rect 62279 -5587 62331 -5577
rect 62139 -5630 62279 -5600
rect 62139 -5640 62140 -5630
rect 61696 -6061 61760 -6059
rect 61888 -6061 61940 -6058
rect 62080 -6061 62140 -5640
rect 62471 -5588 62523 -5578
rect 62331 -5630 62471 -5600
rect 62279 -5649 62331 -5639
rect 62470 -5640 62471 -5630
rect 62661 -5588 62713 -5578
rect 62523 -5630 62661 -5600
rect 62523 -5640 62530 -5630
rect 62470 -6058 62530 -5640
rect 62855 -5588 62907 -5578
rect 62713 -5630 62855 -5600
rect 62661 -5650 62713 -5640
rect 62850 -5640 62855 -5630
rect 63047 -5587 63099 -5577
rect 62907 -5630 63047 -5600
rect 62907 -5640 62910 -5630
rect 62271 -6061 62323 -6059
rect 62464 -6061 62530 -6058
rect 62656 -6061 62708 -6058
rect 62850 -6061 62910 -5640
rect 63238 -5588 63290 -5578
rect 63099 -5630 63238 -5600
rect 63047 -5649 63099 -5639
rect 63230 -5640 63238 -5630
rect 63431 -5588 63483 -5578
rect 63290 -5630 63431 -5600
rect 63041 -6061 63093 -6060
rect 63230 -6061 63290 -5640
rect 63622 -5587 63674 -5577
rect 63483 -5630 63622 -5600
rect 63431 -5650 63483 -5640
rect 63620 -5639 63622 -5630
rect 63814 -5588 63866 -5578
rect 63674 -5630 63814 -5600
rect 63674 -5639 63680 -5630
rect 63620 -6059 63680 -5639
rect 64005 -5588 64057 -5578
rect 63866 -5630 64005 -5600
rect 63814 -5650 63866 -5640
rect 64000 -5640 64005 -5630
rect 64199 -5587 64251 -5577
rect 64057 -5630 64199 -5600
rect 64057 -5640 64060 -5630
rect 64000 -6058 64060 -5640
rect 64390 -5588 64442 -5578
rect 64251 -5630 64390 -5600
rect 64199 -5649 64251 -5639
rect 64582 -5588 64634 -5578
rect 64442 -5630 64582 -5600
rect 64390 -5650 64442 -5640
rect 64774 -5588 64826 -5578
rect 64634 -5630 64774 -5600
rect 64582 -5650 64634 -5640
rect 64966 -5588 65018 -5578
rect 64826 -5630 64966 -5600
rect 64774 -5650 64826 -5640
rect 65159 -5588 65211 -5578
rect 65018 -5630 65159 -5600
rect 64966 -5650 65018 -5640
rect 65350 -5588 65402 -5578
rect 65211 -5630 65350 -5600
rect 65159 -5650 65211 -5640
rect 65543 -5587 65595 -5577
rect 65402 -5630 65543 -5600
rect 65350 -5650 65402 -5640
rect 65734 -5588 65786 -5578
rect 65595 -5630 65734 -5600
rect 65543 -5649 65595 -5639
rect 65927 -5588 65979 -5578
rect 65786 -5630 65927 -5600
rect 65734 -5650 65786 -5640
rect 66118 -5588 66170 -5578
rect 65979 -5630 66118 -5600
rect 65927 -5650 65979 -5640
rect 66309 -5586 66361 -5576
rect 66170 -5630 66309 -5600
rect 66118 -5650 66170 -5640
rect 66504 -5588 66556 -5578
rect 66361 -5630 66504 -5600
rect 66309 -5648 66361 -5638
rect 66504 -5650 66556 -5640
rect 66918 -5950 66970 -5940
rect 66918 -6012 66970 -6002
rect 63423 -6061 63475 -6059
rect 63616 -6061 63680 -6059
rect 63807 -6061 63859 -6058
rect 63998 -6061 64060 -6058
rect 49430 -6074 49482 -6064
rect 49430 -6136 49482 -6126
rect 52047 -6068 64060 -6061
rect 52047 -6069 58623 -6068
rect 52047 -6070 52429 -6069
rect 52047 -6071 52237 -6070
rect 52099 -6092 52237 -6071
rect 52047 -6133 52099 -6123
rect 52289 -6092 52429 -6070
rect 52237 -6132 52289 -6122
rect 52481 -6092 52620 -6069
rect 52429 -6131 52481 -6121
rect 52672 -6092 52814 -6069
rect 52620 -6131 52672 -6121
rect 52866 -6070 53198 -6069
rect 52866 -6092 53004 -6070
rect 52814 -6131 52866 -6121
rect 53056 -6092 53198 -6070
rect 53004 -6132 53056 -6122
rect 53250 -6092 53390 -6069
rect 53198 -6131 53250 -6121
rect 53442 -6070 54542 -6069
rect 53442 -6092 53581 -6070
rect 53390 -6131 53442 -6121
rect 53633 -6092 53776 -6070
rect 53581 -6132 53633 -6122
rect 53828 -6092 53966 -6070
rect 53776 -6132 53828 -6122
rect 54018 -6092 54157 -6070
rect 53966 -6132 54018 -6122
rect 54209 -6092 54349 -6070
rect 54157 -6132 54209 -6122
rect 54401 -6092 54542 -6070
rect 54349 -6132 54401 -6122
rect 54594 -6070 55310 -6069
rect 54594 -6092 54734 -6070
rect 54542 -6131 54594 -6121
rect 54786 -6092 54926 -6070
rect 54734 -6132 54786 -6122
rect 54978 -6092 55119 -6070
rect 54926 -6132 54978 -6122
rect 55171 -6092 55310 -6070
rect 55119 -6132 55171 -6122
rect 55362 -6070 55694 -6069
rect 55362 -6092 55502 -6070
rect 55310 -6131 55362 -6121
rect 55554 -6092 55694 -6070
rect 55502 -6132 55554 -6122
rect 55746 -6092 55886 -6069
rect 55694 -6131 55746 -6121
rect 55938 -6070 56270 -6069
rect 55938 -6092 56077 -6070
rect 55886 -6131 55938 -6121
rect 56129 -6092 56270 -6070
rect 56077 -6132 56129 -6122
rect 56322 -6092 56462 -6069
rect 56270 -6131 56322 -6121
rect 56514 -6070 57613 -6069
rect 56514 -6092 56656 -6070
rect 56462 -6131 56514 -6121
rect 56708 -6071 57036 -6070
rect 56708 -6092 56847 -6071
rect 56656 -6132 56708 -6122
rect 56899 -6092 57036 -6071
rect 56847 -6133 56899 -6123
rect 57088 -6092 57229 -6070
rect 57036 -6132 57088 -6122
rect 57281 -6092 57422 -6070
rect 57229 -6132 57281 -6122
rect 57474 -6092 57613 -6070
rect 57422 -6132 57474 -6122
rect 57665 -6092 57804 -6069
rect 57613 -6131 57665 -6121
rect 57856 -6070 58431 -6069
rect 57856 -6090 58241 -6070
rect 57804 -6131 57856 -6121
rect 58293 -6091 58431 -6070
rect 58241 -6132 58293 -6122
rect 58483 -6091 58623 -6069
rect 58431 -6131 58483 -6121
rect 58675 -6091 58814 -6068
rect 58623 -6130 58675 -6120
rect 58866 -6091 59008 -6068
rect 58814 -6130 58866 -6120
rect 59060 -6069 59392 -6068
rect 59060 -6091 59198 -6069
rect 59008 -6130 59060 -6120
rect 59250 -6091 59392 -6069
rect 59198 -6131 59250 -6121
rect 59444 -6091 59584 -6068
rect 59392 -6130 59444 -6120
rect 59636 -6069 60736 -6068
rect 59636 -6091 59775 -6069
rect 59584 -6130 59636 -6120
rect 59827 -6091 59970 -6069
rect 59775 -6131 59827 -6121
rect 60022 -6091 60160 -6069
rect 59970 -6131 60022 -6121
rect 60212 -6091 60351 -6069
rect 60160 -6131 60212 -6121
rect 60403 -6091 60543 -6069
rect 60351 -6131 60403 -6121
rect 60595 -6091 60736 -6069
rect 60543 -6131 60595 -6121
rect 60788 -6069 61504 -6068
rect 60788 -6091 60928 -6069
rect 60736 -6130 60788 -6120
rect 60980 -6091 61120 -6069
rect 60928 -6131 60980 -6121
rect 61172 -6091 61313 -6069
rect 61120 -6131 61172 -6121
rect 61365 -6091 61504 -6069
rect 61313 -6131 61365 -6121
rect 61556 -6069 61888 -6068
rect 61556 -6091 61696 -6069
rect 61504 -6130 61556 -6120
rect 61748 -6091 61888 -6069
rect 61696 -6131 61748 -6121
rect 61940 -6091 62080 -6068
rect 61888 -6130 61940 -6120
rect 62132 -6069 62464 -6068
rect 62132 -6091 62271 -6069
rect 62080 -6130 62132 -6120
rect 62323 -6091 62464 -6069
rect 62271 -6131 62323 -6121
rect 62516 -6091 62656 -6068
rect 62464 -6130 62516 -6120
rect 62708 -6069 63807 -6068
rect 62708 -6091 62850 -6069
rect 62656 -6130 62708 -6120
rect 62902 -6070 63230 -6069
rect 62902 -6091 63041 -6070
rect 62850 -6131 62902 -6121
rect 63093 -6091 63230 -6070
rect 63041 -6132 63093 -6122
rect 63282 -6091 63423 -6069
rect 63230 -6131 63282 -6121
rect 63475 -6091 63616 -6069
rect 63423 -6131 63475 -6121
rect 63668 -6091 63807 -6069
rect 63616 -6131 63668 -6121
rect 63859 -6091 63998 -6068
rect 63807 -6130 63859 -6120
rect 64050 -6070 64060 -6068
rect 63998 -6130 64050 -6120
rect 49440 -6220 49470 -6136
rect 51949 -6210 52001 -6200
rect 49440 -6260 51949 -6220
rect 47224 -6678 47652 -6264
rect 51116 -6396 51168 -6260
rect 52141 -6210 52193 -6200
rect 52001 -6252 52141 -6222
rect 51949 -6272 52001 -6262
rect 52334 -6210 52386 -6200
rect 52193 -6252 52334 -6222
rect 52141 -6272 52193 -6262
rect 52526 -6210 52578 -6200
rect 52386 -6252 52526 -6222
rect 52334 -6272 52386 -6262
rect 52719 -6210 52771 -6200
rect 52578 -6252 52719 -6222
rect 52526 -6272 52578 -6262
rect 52911 -6209 52963 -6199
rect 52771 -6252 52911 -6222
rect 52719 -6272 52771 -6262
rect 53102 -6210 53154 -6200
rect 52963 -6252 53102 -6222
rect 52911 -6271 52963 -6261
rect 53294 -6210 53346 -6200
rect 53154 -6252 53294 -6222
rect 53102 -6272 53154 -6262
rect 53486 -6209 53538 -6199
rect 53346 -6252 53486 -6222
rect 53294 -6272 53346 -6262
rect 53678 -6209 53730 -6199
rect 53538 -6252 53678 -6222
rect 53486 -6271 53538 -6261
rect 53870 -6210 53922 -6200
rect 53730 -6252 53870 -6222
rect 53678 -6271 53730 -6261
rect 54062 -6209 54114 -6199
rect 53922 -6252 54062 -6222
rect 53870 -6272 53922 -6262
rect 54254 -6210 54306 -6200
rect 54114 -6252 54254 -6222
rect 54062 -6271 54114 -6261
rect 54445 -6209 54497 -6199
rect 54306 -6252 54445 -6222
rect 54254 -6272 54306 -6262
rect 54639 -6210 54691 -6200
rect 54497 -6252 54639 -6222
rect 54445 -6271 54497 -6261
rect 54829 -6210 54881 -6200
rect 54691 -6252 54829 -6222
rect 54639 -6272 54691 -6262
rect 55021 -6210 55073 -6200
rect 54881 -6252 55021 -6222
rect 54829 -6272 54881 -6262
rect 55214 -6210 55266 -6200
rect 55073 -6252 55214 -6222
rect 55021 -6272 55073 -6262
rect 55405 -6210 55457 -6200
rect 55266 -6252 55405 -6222
rect 55214 -6272 55266 -6262
rect 55598 -6209 55650 -6199
rect 55457 -6252 55598 -6222
rect 55405 -6272 55457 -6262
rect 55791 -6210 55843 -6200
rect 55650 -6252 55791 -6222
rect 55598 -6271 55650 -6261
rect 55982 -6210 56034 -6200
rect 55843 -6252 55982 -6222
rect 55791 -6272 55843 -6262
rect 56175 -6210 56227 -6200
rect 56034 -6252 56175 -6222
rect 55982 -6272 56034 -6262
rect 56365 -6210 56417 -6200
rect 56227 -6252 56365 -6222
rect 56175 -6272 56227 -6262
rect 56559 -6209 56611 -6199
rect 56417 -6252 56559 -6222
rect 56365 -6272 56417 -6262
rect 56748 -6210 56800 -6200
rect 56611 -6252 56748 -6222
rect 56559 -6271 56611 -6261
rect 56941 -6210 56993 -6200
rect 56800 -6252 56941 -6222
rect 56748 -6272 56800 -6262
rect 57134 -6210 57186 -6200
rect 56993 -6252 57134 -6222
rect 56941 -6272 56993 -6262
rect 57324 -6210 57376 -6200
rect 57186 -6252 57324 -6222
rect 57134 -6272 57186 -6262
rect 57517 -6209 57569 -6199
rect 57376 -6252 57517 -6222
rect 57324 -6272 57376 -6262
rect 57706 -6209 57758 -6199
rect 57569 -6252 57706 -6222
rect 57517 -6271 57569 -6261
rect 57706 -6271 57758 -6261
rect 58143 -6209 58195 -6199
rect 58335 -6209 58387 -6199
rect 58195 -6251 58335 -6221
rect 58143 -6271 58195 -6261
rect 58528 -6209 58580 -6199
rect 58387 -6251 58528 -6221
rect 58335 -6271 58387 -6261
rect 58720 -6209 58772 -6199
rect 58580 -6251 58720 -6221
rect 58528 -6271 58580 -6261
rect 58913 -6209 58965 -6199
rect 58772 -6251 58913 -6221
rect 58720 -6271 58772 -6261
rect 59105 -6208 59157 -6198
rect 58965 -6251 59105 -6221
rect 58913 -6271 58965 -6261
rect 59296 -6209 59348 -6199
rect 59157 -6251 59296 -6221
rect 59105 -6270 59157 -6260
rect 59488 -6209 59540 -6199
rect 59348 -6251 59488 -6221
rect 59296 -6271 59348 -6261
rect 59680 -6208 59732 -6198
rect 59540 -6251 59680 -6221
rect 59488 -6271 59540 -6261
rect 59872 -6208 59924 -6198
rect 59732 -6251 59872 -6221
rect 59680 -6270 59732 -6260
rect 60064 -6209 60116 -6199
rect 59924 -6251 60064 -6221
rect 59872 -6270 59924 -6260
rect 60256 -6208 60308 -6198
rect 60116 -6251 60256 -6221
rect 60064 -6271 60116 -6261
rect 60448 -6209 60500 -6199
rect 60308 -6251 60448 -6221
rect 60256 -6270 60308 -6260
rect 60639 -6208 60691 -6198
rect 60500 -6251 60639 -6221
rect 60448 -6271 60500 -6261
rect 60833 -6209 60885 -6199
rect 60691 -6251 60833 -6221
rect 60639 -6270 60691 -6260
rect 61023 -6209 61075 -6199
rect 60885 -6251 61023 -6221
rect 60833 -6271 60885 -6261
rect 61215 -6209 61267 -6199
rect 61075 -6251 61215 -6221
rect 61023 -6271 61075 -6261
rect 61408 -6209 61460 -6199
rect 61267 -6251 61408 -6221
rect 61215 -6271 61267 -6261
rect 61599 -6209 61651 -6199
rect 61460 -6251 61599 -6221
rect 61408 -6271 61460 -6261
rect 61792 -6208 61844 -6198
rect 61651 -6251 61792 -6221
rect 61599 -6271 61651 -6261
rect 61985 -6209 62037 -6199
rect 61844 -6251 61985 -6221
rect 61792 -6270 61844 -6260
rect 62176 -6209 62228 -6199
rect 62037 -6251 62176 -6221
rect 61985 -6271 62037 -6261
rect 62369 -6209 62421 -6199
rect 62228 -6251 62369 -6221
rect 62176 -6271 62228 -6261
rect 62559 -6209 62611 -6199
rect 62421 -6251 62559 -6221
rect 62369 -6271 62421 -6261
rect 62753 -6208 62805 -6198
rect 62611 -6251 62753 -6221
rect 62559 -6271 62611 -6261
rect 62942 -6209 62994 -6199
rect 62805 -6251 62942 -6221
rect 62753 -6270 62805 -6260
rect 63135 -6209 63187 -6199
rect 62994 -6251 63135 -6221
rect 62942 -6271 62994 -6261
rect 63328 -6209 63380 -6199
rect 63187 -6251 63328 -6221
rect 63135 -6271 63187 -6261
rect 63518 -6209 63570 -6199
rect 63380 -6251 63518 -6221
rect 63328 -6271 63380 -6261
rect 63711 -6208 63763 -6198
rect 63570 -6251 63711 -6221
rect 63518 -6271 63570 -6261
rect 63900 -6208 63952 -6198
rect 63763 -6251 63900 -6221
rect 63711 -6270 63763 -6260
rect 66930 -6220 66960 -6012
rect 63952 -6250 66960 -6220
rect 63900 -6270 63952 -6260
rect 63990 -6300 64050 -6290
rect 57800 -6310 57860 -6300
rect 51116 -6458 51168 -6448
rect 52040 -6320 52100 -6310
rect 47224 -7752 47254 -6678
rect 47614 -7752 47652 -6678
rect 51116 -6500 51168 -6490
rect 51116 -6680 51168 -6552
rect 52040 -6680 52100 -6380
rect 52238 -6680 52290 -6678
rect 52430 -6680 52482 -6677
rect 52621 -6680 52673 -6677
rect 52815 -6680 52867 -6677
rect 53005 -6680 53057 -6678
rect 53199 -6680 53251 -6677
rect 53391 -6680 53443 -6677
rect 53582 -6680 53634 -6678
rect 53777 -6680 53829 -6678
rect 53967 -6680 54019 -6678
rect 54158 -6680 54210 -6678
rect 54350 -6680 54402 -6678
rect 54543 -6680 54595 -6677
rect 54735 -6680 54787 -6678
rect 54927 -6680 54979 -6678
rect 55120 -6680 55172 -6678
rect 55311 -6680 55363 -6677
rect 55503 -6680 55555 -6678
rect 55695 -6680 55747 -6677
rect 55887 -6680 55939 -6677
rect 56078 -6680 56130 -6678
rect 56271 -6680 56323 -6677
rect 56463 -6680 56515 -6677
rect 56657 -6680 56709 -6678
rect 56848 -6680 56900 -6679
rect 57037 -6680 57089 -6678
rect 57230 -6680 57282 -6678
rect 57423 -6680 57475 -6678
rect 57614 -6680 57666 -6677
rect 57800 -6680 57860 -6370
rect 49440 -6687 57860 -6680
rect 49440 -6688 52430 -6687
rect 49440 -6689 52238 -6688
rect 49440 -6720 52048 -6689
rect 49440 -6862 49470 -6720
rect 52100 -6710 52238 -6689
rect 52048 -6751 52100 -6741
rect 52290 -6710 52430 -6688
rect 52238 -6750 52290 -6740
rect 52482 -6710 52621 -6687
rect 52430 -6749 52482 -6739
rect 52673 -6710 52815 -6687
rect 52621 -6749 52673 -6739
rect 52867 -6688 53199 -6687
rect 52867 -6710 53005 -6688
rect 52815 -6749 52867 -6739
rect 53057 -6710 53199 -6688
rect 53005 -6750 53057 -6740
rect 53251 -6710 53391 -6687
rect 53199 -6749 53251 -6739
rect 53443 -6688 54543 -6687
rect 53443 -6710 53582 -6688
rect 53391 -6749 53443 -6739
rect 53634 -6710 53777 -6688
rect 53582 -6750 53634 -6740
rect 53829 -6710 53967 -6688
rect 53777 -6750 53829 -6740
rect 54019 -6710 54158 -6688
rect 53967 -6750 54019 -6740
rect 54210 -6710 54350 -6688
rect 54158 -6750 54210 -6740
rect 54402 -6710 54543 -6688
rect 54350 -6750 54402 -6740
rect 54595 -6688 55311 -6687
rect 54595 -6710 54735 -6688
rect 54543 -6749 54595 -6739
rect 54787 -6710 54927 -6688
rect 54735 -6750 54787 -6740
rect 54979 -6710 55120 -6688
rect 54927 -6750 54979 -6740
rect 55172 -6710 55311 -6688
rect 55120 -6750 55172 -6740
rect 55363 -6688 55695 -6687
rect 55363 -6710 55503 -6688
rect 55311 -6749 55363 -6739
rect 55555 -6710 55695 -6688
rect 55503 -6750 55555 -6740
rect 55747 -6710 55887 -6687
rect 55695 -6749 55747 -6739
rect 55939 -6688 56271 -6687
rect 55939 -6710 56078 -6688
rect 55887 -6749 55939 -6739
rect 56130 -6710 56271 -6688
rect 56078 -6750 56130 -6740
rect 56323 -6710 56463 -6687
rect 56271 -6749 56323 -6739
rect 56515 -6688 57614 -6687
rect 56515 -6710 56657 -6688
rect 56463 -6749 56515 -6739
rect 56709 -6689 57037 -6688
rect 56709 -6710 56848 -6689
rect 56657 -6750 56709 -6740
rect 56900 -6710 57037 -6689
rect 56848 -6751 56900 -6741
rect 57089 -6710 57230 -6688
rect 57037 -6750 57089 -6740
rect 57282 -6710 57423 -6688
rect 57230 -6750 57282 -6740
rect 57475 -6710 57614 -6688
rect 57423 -6750 57475 -6740
rect 57666 -6710 57805 -6687
rect 57614 -6749 57666 -6739
rect 57857 -6690 57860 -6687
rect 58230 -6310 58290 -6300
rect 58230 -6679 58290 -6370
rect 58426 -6679 58478 -6677
rect 58618 -6679 58670 -6676
rect 58809 -6679 58861 -6676
rect 59003 -6679 59055 -6676
rect 59193 -6679 59245 -6677
rect 59387 -6679 59439 -6676
rect 59579 -6679 59631 -6676
rect 59770 -6679 59822 -6677
rect 59965 -6679 60017 -6677
rect 60155 -6679 60207 -6677
rect 60346 -6679 60398 -6677
rect 60538 -6679 60590 -6677
rect 60731 -6679 60783 -6676
rect 60923 -6679 60975 -6677
rect 61115 -6679 61167 -6677
rect 61308 -6679 61360 -6677
rect 61499 -6679 61551 -6676
rect 61691 -6679 61743 -6677
rect 61883 -6679 61935 -6676
rect 62075 -6679 62127 -6676
rect 62266 -6679 62318 -6677
rect 62459 -6679 62511 -6676
rect 62651 -6679 62703 -6676
rect 62845 -6679 62897 -6677
rect 63036 -6679 63088 -6678
rect 63225 -6679 63277 -6677
rect 63418 -6679 63470 -6677
rect 63611 -6679 63663 -6677
rect 63802 -6679 63854 -6676
rect 63990 -6679 64050 -6360
rect 64530 -6380 64582 -6250
rect 64530 -6442 64582 -6432
rect 68894 -6272 68930 -5188
rect 69296 -6272 69326 -5188
rect 58230 -6680 64050 -6679
rect 64536 -6496 64588 -6486
rect 64536 -6680 64588 -6548
rect 68894 -6672 69326 -6272
rect 58230 -6686 66950 -6680
rect 58230 -6687 58618 -6686
rect 58230 -6688 58426 -6687
rect 58230 -6690 58236 -6688
rect 57805 -6749 57857 -6739
rect 58288 -6709 58426 -6688
rect 58236 -6750 58288 -6740
rect 58478 -6709 58618 -6687
rect 58426 -6749 58478 -6739
rect 58670 -6709 58809 -6686
rect 58618 -6748 58670 -6738
rect 58861 -6709 59003 -6686
rect 58809 -6748 58861 -6738
rect 59055 -6687 59387 -6686
rect 59055 -6709 59193 -6687
rect 59003 -6748 59055 -6738
rect 59245 -6709 59387 -6687
rect 59193 -6749 59245 -6739
rect 59439 -6709 59579 -6686
rect 59387 -6748 59439 -6738
rect 59631 -6687 60731 -6686
rect 59631 -6709 59770 -6687
rect 59579 -6748 59631 -6738
rect 59822 -6709 59965 -6687
rect 59770 -6749 59822 -6739
rect 60017 -6709 60155 -6687
rect 59965 -6749 60017 -6739
rect 60207 -6709 60346 -6687
rect 60155 -6749 60207 -6739
rect 60398 -6709 60538 -6687
rect 60346 -6749 60398 -6739
rect 60590 -6709 60731 -6687
rect 60538 -6749 60590 -6739
rect 60783 -6687 61499 -6686
rect 60783 -6709 60923 -6687
rect 60731 -6748 60783 -6738
rect 60975 -6709 61115 -6687
rect 60923 -6749 60975 -6739
rect 61167 -6709 61308 -6687
rect 61115 -6749 61167 -6739
rect 61360 -6709 61499 -6687
rect 61308 -6749 61360 -6739
rect 61551 -6687 61883 -6686
rect 61551 -6709 61691 -6687
rect 61499 -6748 61551 -6738
rect 61743 -6709 61883 -6687
rect 61691 -6749 61743 -6739
rect 61935 -6709 62075 -6686
rect 61883 -6748 61935 -6738
rect 62127 -6687 62459 -6686
rect 62127 -6709 62266 -6687
rect 62075 -6748 62127 -6738
rect 62318 -6709 62459 -6687
rect 62266 -6749 62318 -6739
rect 62511 -6709 62651 -6686
rect 62459 -6748 62511 -6738
rect 62703 -6687 63802 -6686
rect 62703 -6709 62845 -6687
rect 62651 -6748 62703 -6738
rect 62897 -6688 63225 -6687
rect 62897 -6709 63036 -6688
rect 62845 -6749 62897 -6739
rect 63088 -6709 63225 -6688
rect 63036 -6750 63088 -6740
rect 63277 -6709 63418 -6687
rect 63225 -6749 63277 -6739
rect 63470 -6709 63611 -6687
rect 63418 -6749 63470 -6739
rect 63663 -6709 63802 -6687
rect 63611 -6749 63663 -6739
rect 63854 -6709 63993 -6686
rect 63802 -6748 63854 -6738
rect 64045 -6710 66950 -6686
rect 63993 -6748 64045 -6738
rect 51950 -6826 63950 -6810
rect 51950 -6827 59100 -6826
rect 51950 -6828 52912 -6827
rect 49436 -6872 49488 -6862
rect 52002 -6880 52142 -6828
rect 52194 -6880 52335 -6828
rect 52387 -6880 52527 -6828
rect 52579 -6880 52720 -6828
rect 52772 -6879 52912 -6828
rect 52964 -6828 53487 -6827
rect 52964 -6879 53103 -6828
rect 52772 -6880 53103 -6879
rect 53155 -6880 53295 -6828
rect 53347 -6879 53487 -6828
rect 53539 -6879 53679 -6827
rect 53731 -6828 54063 -6827
rect 53731 -6879 53871 -6828
rect 53347 -6880 53871 -6879
rect 53923 -6879 54063 -6828
rect 54115 -6828 54446 -6827
rect 54115 -6879 54255 -6828
rect 53923 -6880 54255 -6879
rect 54307 -6879 54446 -6828
rect 54498 -6828 55599 -6827
rect 54498 -6879 54640 -6828
rect 54307 -6880 54640 -6879
rect 54692 -6880 54830 -6828
rect 54882 -6880 55022 -6828
rect 55074 -6880 55215 -6828
rect 55267 -6880 55406 -6828
rect 55458 -6879 55599 -6828
rect 55651 -6828 56560 -6827
rect 55651 -6879 55792 -6828
rect 55458 -6880 55792 -6879
rect 55844 -6880 55983 -6828
rect 56035 -6880 56176 -6828
rect 56228 -6880 56366 -6828
rect 56418 -6879 56560 -6828
rect 56612 -6828 57518 -6827
rect 56612 -6879 56749 -6828
rect 56418 -6880 56749 -6879
rect 56801 -6880 56942 -6828
rect 56994 -6880 57135 -6828
rect 57187 -6880 57325 -6828
rect 57377 -6879 57518 -6828
rect 57570 -6879 57707 -6827
rect 57759 -6879 58138 -6827
rect 58190 -6879 58330 -6827
rect 58382 -6879 58523 -6827
rect 58575 -6879 58715 -6827
rect 58767 -6879 58908 -6827
rect 58960 -6878 59100 -6827
rect 59152 -6827 59675 -6826
rect 59152 -6878 59291 -6827
rect 58960 -6879 59291 -6878
rect 59343 -6879 59483 -6827
rect 59535 -6878 59675 -6827
rect 59727 -6878 59867 -6826
rect 59919 -6827 60251 -6826
rect 59919 -6878 60059 -6827
rect 59535 -6879 60059 -6878
rect 60111 -6878 60251 -6827
rect 60303 -6827 60634 -6826
rect 60303 -6878 60443 -6827
rect 60111 -6879 60443 -6878
rect 60495 -6878 60634 -6827
rect 60686 -6827 61787 -6826
rect 60686 -6878 60828 -6827
rect 60495 -6879 60828 -6878
rect 60880 -6879 61018 -6827
rect 61070 -6879 61210 -6827
rect 61262 -6879 61403 -6827
rect 61455 -6879 61594 -6827
rect 61646 -6878 61787 -6827
rect 61839 -6827 62748 -6826
rect 61839 -6878 61980 -6827
rect 61646 -6879 61980 -6878
rect 62032 -6879 62171 -6827
rect 62223 -6879 62364 -6827
rect 62416 -6879 62554 -6827
rect 62606 -6878 62748 -6827
rect 62800 -6827 63706 -6826
rect 62800 -6878 62937 -6827
rect 62606 -6879 62937 -6878
rect 62989 -6879 63130 -6827
rect 63182 -6879 63323 -6827
rect 63375 -6879 63513 -6827
rect 63565 -6878 63706 -6827
rect 63758 -6878 63895 -6826
rect 63947 -6878 63950 -6826
rect 66920 -6840 66950 -6710
rect 63565 -6879 63950 -6878
rect 57377 -6880 63950 -6879
rect 51950 -6890 63950 -6880
rect 66912 -6850 66964 -6840
rect 49436 -6934 49488 -6924
rect 50087 -7300 50139 -7292
rect 50277 -7300 50329 -7291
rect 50470 -7300 50522 -7294
rect 50662 -7299 50714 -7289
rect 50087 -7301 50662 -7300
rect 50087 -7302 50277 -7301
rect 50139 -7330 50277 -7302
rect 50087 -7364 50139 -7354
rect 50329 -7304 50662 -7301
rect 50329 -7330 50470 -7304
rect 50277 -7363 50329 -7353
rect 50522 -7330 50662 -7304
rect 50470 -7366 50522 -7356
rect 50854 -7300 50906 -7293
rect 51046 -7298 51098 -7288
rect 50714 -7303 51046 -7300
rect 50714 -7330 50854 -7303
rect 50662 -7361 50714 -7351
rect 50906 -7330 51046 -7303
rect 50854 -7365 50906 -7355
rect 51238 -7299 51290 -7289
rect 51098 -7330 51238 -7300
rect 51046 -7360 51098 -7350
rect 51428 -7298 51480 -7288
rect 51290 -7330 51428 -7300
rect 51238 -7361 51290 -7351
rect 51622 -7300 51674 -7299
rect 51811 -7300 51863 -7297
rect 52000 -7300 52060 -6890
rect 52200 -7300 52252 -7298
rect 52390 -7300 52450 -6890
rect 52582 -7300 52634 -7298
rect 52774 -7300 52826 -7291
rect 52960 -7300 53020 -6890
rect 53159 -7300 53211 -7292
rect 53350 -7300 53410 -6890
rect 53542 -7300 53594 -7290
rect 53730 -7300 53790 -6890
rect 54120 -7287 54180 -6890
rect 53927 -7300 53979 -7291
rect 54119 -7297 54180 -7287
rect 54510 -7291 54570 -6890
rect 54890 -7290 54950 -6890
rect 55260 -7288 55320 -6890
rect 51480 -7301 53351 -7300
rect 51480 -7307 52774 -7301
rect 51480 -7309 51811 -7307
rect 51480 -7330 51622 -7309
rect 51428 -7360 51480 -7350
rect 51674 -7330 51811 -7309
rect 51622 -7371 51674 -7361
rect 51863 -7330 52001 -7307
rect 51811 -7369 51863 -7359
rect 52053 -7308 52392 -7307
rect 52053 -7330 52200 -7308
rect 52001 -7369 52053 -7359
rect 52252 -7330 52392 -7308
rect 52200 -7370 52252 -7360
rect 52444 -7308 52774 -7307
rect 52444 -7330 52582 -7308
rect 52392 -7369 52444 -7359
rect 52634 -7330 52774 -7308
rect 52582 -7370 52634 -7360
rect 52826 -7302 53351 -7301
rect 52826 -7303 53159 -7302
rect 52826 -7330 52966 -7303
rect 52774 -7363 52826 -7353
rect 53018 -7330 53159 -7303
rect 52966 -7365 53018 -7355
rect 53211 -7330 53351 -7302
rect 53159 -7364 53211 -7354
rect 53403 -7330 53542 -7300
rect 53351 -7362 53403 -7352
rect 53594 -7301 54119 -7300
rect 53594 -7305 53927 -7301
rect 53594 -7330 53736 -7305
rect 53542 -7362 53594 -7352
rect 53788 -7330 53927 -7305
rect 53736 -7367 53788 -7357
rect 53979 -7330 54119 -7301
rect 53927 -7363 53979 -7353
rect 54171 -7300 54180 -7297
rect 54312 -7300 54364 -7291
rect 54504 -7300 54570 -7291
rect 54697 -7300 54749 -7292
rect 54889 -7300 54950 -7290
rect 55080 -7299 55132 -7289
rect 54171 -7301 54889 -7300
rect 54171 -7330 54312 -7301
rect 54119 -7359 54171 -7349
rect 54364 -7330 54504 -7301
rect 54312 -7363 54364 -7353
rect 54556 -7302 54889 -7301
rect 54556 -7330 54697 -7302
rect 54504 -7363 54556 -7353
rect 54749 -7330 54889 -7302
rect 54697 -7364 54749 -7354
rect 54941 -7330 55080 -7300
rect 54889 -7362 54941 -7352
rect 55260 -7298 55323 -7288
rect 55260 -7300 55271 -7298
rect 55132 -7330 55271 -7300
rect 55080 -7361 55132 -7351
rect 55464 -7298 55516 -7288
rect 55323 -7330 55464 -7300
rect 55271 -7360 55323 -7350
rect 55650 -7300 55710 -6890
rect 55846 -7300 55898 -7298
rect 56030 -7300 56090 -6890
rect 56410 -7300 56470 -6890
rect 56810 -7300 56870 -6890
rect 57180 -7296 57240 -6890
rect 56997 -7300 57049 -7298
rect 57180 -7300 57243 -7296
rect 57384 -7300 57436 -7297
rect 57570 -7300 57630 -6890
rect 57960 -7298 58020 -6890
rect 57766 -7300 57818 -7298
rect 57959 -7300 58020 -7298
rect 58151 -7300 58203 -7298
rect 58340 -7300 58400 -6890
rect 58730 -7297 58790 -6890
rect 58535 -7300 58587 -7298
rect 58726 -7300 58790 -7297
rect 58921 -7300 58973 -7298
rect 59110 -7300 59170 -6890
rect 59303 -7300 59355 -7298
rect 59490 -7300 59550 -6890
rect 59880 -7298 59940 -6890
rect 59686 -7300 59738 -7298
rect 59878 -7300 59940 -7298
rect 60071 -7300 60123 -7298
rect 60260 -7300 60320 -6890
rect 60454 -7300 60506 -7298
rect 60640 -7300 60700 -6890
rect 60838 -7300 60890 -7298
rect 61030 -7300 61090 -6890
rect 61420 -7297 61480 -6890
rect 61222 -7300 61274 -7299
rect 61415 -7300 61480 -7297
rect 61605 -7300 61657 -7297
rect 61800 -7299 61860 -6890
rect 61798 -7300 61860 -7299
rect 61990 -7300 62042 -7298
rect 62180 -7300 62240 -6890
rect 62374 -7300 62426 -7297
rect 62570 -7298 62630 -6890
rect 62950 -7298 63010 -6890
rect 62566 -7300 62630 -7298
rect 62757 -7300 62809 -7298
rect 62949 -7300 63010 -7298
rect 63143 -7300 63195 -7297
rect 63340 -7298 63400 -6890
rect 63335 -7300 63400 -7298
rect 63525 -7300 63577 -7299
rect 63720 -7300 63780 -6890
rect 66912 -6912 66964 -6902
rect 63909 -7300 63961 -7298
rect 64102 -7300 64154 -7297
rect 64295 -7300 64347 -7298
rect 64486 -7300 64538 -7298
rect 64677 -7300 64729 -7298
rect 64870 -7300 64922 -7298
rect 65063 -7300 65115 -7298
rect 65254 -7300 65306 -7298
rect 65445 -7300 65497 -7297
rect 65636 -7300 65688 -7297
rect 65829 -7300 65881 -7298
rect 66023 -7300 66075 -7298
rect 66211 -7300 66263 -7299
rect 55516 -7306 66470 -7300
rect 55516 -7307 57191 -7306
rect 55516 -7330 55655 -7307
rect 55464 -7360 55516 -7350
rect 55707 -7308 57191 -7307
rect 55707 -7330 55846 -7308
rect 55655 -7369 55707 -7359
rect 55898 -7309 56997 -7308
rect 55898 -7330 56036 -7309
rect 55846 -7370 55898 -7360
rect 56088 -7311 56997 -7309
rect 56088 -7313 56808 -7311
rect 56088 -7330 56230 -7313
rect 56036 -7371 56088 -7361
rect 56282 -7314 56808 -7313
rect 56282 -7315 56616 -7314
rect 56282 -7330 56422 -7315
rect 56230 -7375 56282 -7365
rect 56474 -7330 56616 -7315
rect 56422 -7377 56474 -7367
rect 56668 -7330 56808 -7314
rect 56616 -7376 56668 -7366
rect 56860 -7330 56997 -7311
rect 56808 -7373 56860 -7363
rect 57049 -7330 57191 -7308
rect 56997 -7370 57049 -7360
rect 57243 -7307 66470 -7306
rect 57243 -7330 57384 -7307
rect 57191 -7368 57243 -7358
rect 57436 -7308 58726 -7307
rect 57436 -7330 57577 -7308
rect 57384 -7369 57436 -7359
rect 57629 -7330 57766 -7308
rect 57577 -7370 57629 -7360
rect 57818 -7330 57959 -7308
rect 57766 -7370 57818 -7360
rect 58011 -7330 58151 -7308
rect 57959 -7370 58011 -7360
rect 58203 -7330 58342 -7308
rect 58151 -7370 58203 -7360
rect 58394 -7330 58535 -7308
rect 58342 -7370 58394 -7360
rect 58587 -7330 58726 -7308
rect 58535 -7370 58587 -7360
rect 58778 -7308 61415 -7307
rect 58778 -7330 58921 -7308
rect 58726 -7369 58778 -7359
rect 58973 -7330 59110 -7308
rect 58921 -7370 58973 -7360
rect 59162 -7330 59303 -7308
rect 59110 -7370 59162 -7360
rect 59355 -7330 59495 -7308
rect 59303 -7370 59355 -7360
rect 59547 -7330 59686 -7308
rect 59495 -7370 59547 -7360
rect 59738 -7330 59878 -7308
rect 59686 -7370 59738 -7360
rect 59930 -7330 60071 -7308
rect 59878 -7370 59930 -7360
rect 60123 -7309 60454 -7308
rect 60123 -7330 60260 -7309
rect 60071 -7370 60123 -7360
rect 60312 -7330 60454 -7309
rect 60260 -7371 60312 -7361
rect 60506 -7330 60645 -7308
rect 60454 -7370 60506 -7360
rect 60697 -7330 60838 -7308
rect 60645 -7370 60697 -7360
rect 60890 -7330 61030 -7308
rect 60838 -7370 60890 -7360
rect 61082 -7309 61415 -7308
rect 61082 -7330 61222 -7309
rect 61030 -7370 61082 -7360
rect 61274 -7330 61415 -7309
rect 61222 -7371 61274 -7361
rect 61467 -7330 61605 -7307
rect 61415 -7369 61467 -7359
rect 61657 -7308 62183 -7307
rect 61657 -7309 61990 -7308
rect 61657 -7330 61798 -7309
rect 61605 -7369 61657 -7359
rect 61850 -7330 61990 -7309
rect 61798 -7371 61850 -7361
rect 62042 -7330 62183 -7308
rect 61990 -7370 62042 -7360
rect 62235 -7330 62374 -7307
rect 62183 -7369 62235 -7359
rect 62426 -7308 63143 -7307
rect 62426 -7330 62566 -7308
rect 62374 -7369 62426 -7359
rect 62618 -7330 62757 -7308
rect 62566 -7370 62618 -7360
rect 62809 -7330 62949 -7308
rect 62757 -7370 62809 -7360
rect 63001 -7330 63143 -7308
rect 62949 -7370 63001 -7360
rect 63195 -7308 64102 -7307
rect 63195 -7330 63335 -7308
rect 63143 -7369 63195 -7359
rect 63387 -7309 63909 -7308
rect 63387 -7330 63525 -7309
rect 63335 -7370 63387 -7360
rect 63577 -7310 63909 -7309
rect 63577 -7330 63716 -7310
rect 63525 -7371 63577 -7361
rect 63768 -7330 63909 -7310
rect 63716 -7372 63768 -7362
rect 63961 -7330 64102 -7308
rect 63909 -7370 63961 -7360
rect 64154 -7308 65445 -7307
rect 64154 -7330 64295 -7308
rect 64102 -7369 64154 -7359
rect 64347 -7330 64486 -7308
rect 64295 -7370 64347 -7360
rect 64538 -7330 64677 -7308
rect 64486 -7370 64538 -7360
rect 64729 -7330 64870 -7308
rect 64677 -7370 64729 -7360
rect 64922 -7330 65063 -7308
rect 64870 -7370 64922 -7360
rect 65115 -7330 65254 -7308
rect 65063 -7370 65115 -7360
rect 65306 -7330 65445 -7308
rect 65254 -7370 65306 -7360
rect 65497 -7330 65636 -7307
rect 65445 -7369 65497 -7359
rect 65688 -7308 66470 -7307
rect 65688 -7330 65829 -7308
rect 65636 -7369 65688 -7359
rect 65881 -7330 66023 -7308
rect 65829 -7370 65881 -7360
rect 66075 -7309 66470 -7308
rect 66075 -7330 66211 -7309
rect 66023 -7370 66075 -7360
rect 66263 -7317 66470 -7309
rect 66263 -7330 66405 -7317
rect 66211 -7371 66263 -7361
rect 66457 -7330 66470 -7317
rect 66405 -7379 66457 -7369
rect 49991 -7445 50043 -7435
rect 50182 -7447 50234 -7437
rect 50043 -7490 50182 -7460
rect 50043 -7497 50070 -7490
rect 49991 -7507 50070 -7497
rect 50000 -7654 50070 -7507
rect 50374 -7446 50426 -7436
rect 50234 -7490 50374 -7460
rect 50182 -7509 50234 -7499
rect 50566 -7449 50618 -7439
rect 50426 -7490 50566 -7460
rect 50374 -7508 50426 -7498
rect 50760 -7448 50812 -7438
rect 50618 -7490 50760 -7460
rect 50566 -7511 50618 -7501
rect 50950 -7448 51002 -7438
rect 50812 -7490 50950 -7460
rect 50760 -7510 50812 -7500
rect 51145 -7446 51197 -7436
rect 51002 -7490 51145 -7460
rect 50950 -7510 51002 -7500
rect 51336 -7445 51388 -7435
rect 51197 -7490 51336 -7460
rect 51145 -7508 51197 -7498
rect 51531 -7447 51583 -7437
rect 51388 -7490 51531 -7460
rect 51336 -7507 51388 -7497
rect 51721 -7447 51773 -7437
rect 51583 -7490 51721 -7460
rect 51531 -7509 51583 -7499
rect 51911 -7446 51963 -7436
rect 51773 -7490 51911 -7460
rect 51721 -7509 51773 -7499
rect 52104 -7445 52156 -7435
rect 51963 -7490 52104 -7460
rect 51911 -7508 51963 -7498
rect 52295 -7445 52347 -7435
rect 52156 -7490 52295 -7460
rect 52104 -7507 52156 -7497
rect 52491 -7447 52543 -7437
rect 52347 -7490 52491 -7460
rect 52295 -7507 52347 -7497
rect 52680 -7447 52732 -7437
rect 52543 -7490 52680 -7460
rect 52491 -7509 52543 -7499
rect 52874 -7447 52926 -7437
rect 52732 -7490 52874 -7460
rect 52680 -7509 52732 -7499
rect 53063 -7447 53115 -7437
rect 52926 -7490 53063 -7460
rect 52874 -7509 52926 -7499
rect 53255 -7448 53307 -7438
rect 53115 -7490 53255 -7460
rect 53063 -7509 53115 -7499
rect 53448 -7448 53500 -7438
rect 53307 -7490 53448 -7460
rect 53255 -7510 53307 -7500
rect 53639 -7448 53691 -7438
rect 53500 -7490 53639 -7460
rect 53448 -7510 53500 -7500
rect 53831 -7447 53883 -7437
rect 53691 -7490 53831 -7460
rect 53639 -7510 53691 -7500
rect 54023 -7448 54075 -7438
rect 53883 -7490 54023 -7460
rect 53831 -7509 53883 -7499
rect 54216 -7448 54268 -7438
rect 54075 -7490 54216 -7460
rect 54023 -7510 54075 -7500
rect 54407 -7448 54459 -7438
rect 54268 -7490 54407 -7460
rect 54216 -7510 54268 -7500
rect 54599 -7447 54651 -7437
rect 54459 -7490 54599 -7460
rect 54407 -7510 54459 -7500
rect 54792 -7448 54844 -7438
rect 54651 -7490 54792 -7460
rect 54599 -7509 54651 -7499
rect 54984 -7448 55036 -7438
rect 54844 -7490 54984 -7460
rect 54792 -7510 54844 -7500
rect 55175 -7448 55227 -7438
rect 55036 -7490 55175 -7460
rect 54984 -7510 55036 -7500
rect 55366 -7448 55418 -7438
rect 55227 -7490 55366 -7460
rect 55175 -7510 55227 -7500
rect 55558 -7448 55610 -7438
rect 55418 -7490 55558 -7460
rect 55366 -7510 55418 -7500
rect 55751 -7447 55803 -7437
rect 55610 -7490 55751 -7460
rect 55558 -7510 55610 -7500
rect 55942 -7447 55994 -7437
rect 55803 -7490 55942 -7460
rect 55751 -7509 55803 -7499
rect 56136 -7448 56188 -7438
rect 55994 -7490 56136 -7460
rect 55942 -7509 55994 -7499
rect 56328 -7448 56380 -7438
rect 56188 -7490 56328 -7460
rect 56136 -7510 56188 -7500
rect 56520 -7448 56572 -7438
rect 56380 -7490 56520 -7460
rect 56328 -7510 56380 -7500
rect 56712 -7448 56764 -7438
rect 56572 -7490 56712 -7460
rect 56520 -7510 56572 -7500
rect 56904 -7448 56956 -7438
rect 56764 -7490 56904 -7460
rect 56712 -7510 56764 -7500
rect 57096 -7448 57148 -7438
rect 56956 -7490 57096 -7460
rect 56904 -7510 56956 -7500
rect 57288 -7448 57340 -7438
rect 57148 -7490 57288 -7460
rect 57096 -7510 57148 -7500
rect 57479 -7448 57531 -7438
rect 57340 -7490 57479 -7460
rect 57288 -7510 57340 -7500
rect 57671 -7448 57723 -7438
rect 57531 -7490 57671 -7460
rect 57479 -7510 57531 -7500
rect 57864 -7448 57916 -7438
rect 57723 -7490 57864 -7460
rect 57671 -7510 57723 -7500
rect 58056 -7448 58108 -7438
rect 57916 -7490 58056 -7460
rect 57864 -7510 57916 -7500
rect 58248 -7448 58300 -7438
rect 58108 -7490 58248 -7460
rect 58056 -7510 58108 -7500
rect 58439 -7448 58491 -7438
rect 58300 -7490 58439 -7460
rect 58248 -7510 58300 -7500
rect 58631 -7448 58683 -7438
rect 58491 -7490 58631 -7460
rect 58439 -7510 58491 -7500
rect 58822 -7448 58874 -7438
rect 58683 -7490 58822 -7460
rect 58631 -7510 58683 -7500
rect 59013 -7448 59065 -7438
rect 58874 -7490 59013 -7460
rect 58822 -7510 58874 -7500
rect 59207 -7448 59259 -7438
rect 59065 -7490 59207 -7460
rect 59013 -7510 59065 -7500
rect 59399 -7448 59451 -7438
rect 59259 -7490 59399 -7460
rect 59207 -7510 59259 -7500
rect 59592 -7447 59644 -7437
rect 59451 -7490 59592 -7460
rect 59399 -7510 59451 -7500
rect 59783 -7448 59835 -7438
rect 59644 -7490 59783 -7460
rect 59592 -7509 59644 -7499
rect 59975 -7448 60027 -7438
rect 59835 -7490 59975 -7460
rect 59783 -7510 59835 -7500
rect 60168 -7448 60220 -7438
rect 60027 -7490 60168 -7460
rect 59975 -7510 60027 -7500
rect 60360 -7448 60412 -7438
rect 60220 -7490 60360 -7460
rect 60168 -7510 60220 -7500
rect 60553 -7447 60605 -7437
rect 60412 -7490 60553 -7460
rect 60360 -7510 60412 -7500
rect 60744 -7448 60796 -7438
rect 60605 -7490 60744 -7460
rect 60553 -7509 60605 -7499
rect 60936 -7448 60988 -7438
rect 60796 -7490 60936 -7460
rect 60744 -7510 60796 -7500
rect 61127 -7448 61179 -7438
rect 60988 -7490 61127 -7460
rect 60936 -7510 60988 -7500
rect 61319 -7448 61371 -7438
rect 61179 -7490 61319 -7460
rect 61127 -7510 61179 -7500
rect 61511 -7448 61563 -7438
rect 61371 -7490 61511 -7460
rect 61319 -7510 61371 -7500
rect 61704 -7448 61756 -7438
rect 61563 -7490 61704 -7460
rect 61511 -7510 61563 -7500
rect 61895 -7448 61947 -7438
rect 61756 -7490 61895 -7460
rect 61704 -7510 61756 -7500
rect 62087 -7448 62139 -7438
rect 61947 -7490 62087 -7460
rect 61895 -7510 61947 -7500
rect 62279 -7447 62331 -7437
rect 62139 -7490 62279 -7460
rect 62087 -7510 62139 -7500
rect 62471 -7448 62523 -7438
rect 62331 -7490 62471 -7460
rect 62279 -7509 62331 -7499
rect 62661 -7448 62713 -7438
rect 62523 -7490 62661 -7460
rect 62471 -7510 62523 -7500
rect 62855 -7448 62907 -7438
rect 62713 -7490 62855 -7460
rect 62661 -7510 62713 -7500
rect 63047 -7447 63099 -7437
rect 62907 -7490 63047 -7460
rect 62855 -7510 62907 -7500
rect 63238 -7448 63290 -7438
rect 63099 -7490 63238 -7460
rect 63047 -7509 63099 -7499
rect 63431 -7448 63483 -7438
rect 63290 -7490 63431 -7460
rect 63238 -7510 63290 -7500
rect 63622 -7447 63674 -7437
rect 63483 -7490 63622 -7460
rect 63431 -7510 63483 -7500
rect 63814 -7448 63866 -7438
rect 63674 -7490 63814 -7460
rect 63622 -7509 63674 -7499
rect 64005 -7448 64057 -7438
rect 63866 -7490 64005 -7460
rect 63814 -7510 63866 -7500
rect 64199 -7447 64251 -7437
rect 64057 -7490 64199 -7460
rect 64005 -7510 64057 -7500
rect 64390 -7448 64442 -7438
rect 64251 -7490 64390 -7460
rect 64199 -7509 64251 -7499
rect 64582 -7448 64634 -7438
rect 64442 -7490 64582 -7460
rect 64390 -7510 64442 -7500
rect 64774 -7448 64826 -7438
rect 64634 -7490 64774 -7460
rect 64582 -7510 64634 -7500
rect 64966 -7448 65018 -7438
rect 64826 -7490 64966 -7460
rect 64774 -7510 64826 -7500
rect 65159 -7448 65211 -7438
rect 65018 -7490 65159 -7460
rect 64966 -7510 65018 -7500
rect 65350 -7448 65402 -7438
rect 65211 -7490 65350 -7460
rect 65159 -7510 65211 -7500
rect 65543 -7447 65595 -7437
rect 65402 -7490 65543 -7460
rect 65350 -7510 65402 -7500
rect 65734 -7448 65786 -7438
rect 65595 -7490 65734 -7460
rect 65543 -7509 65595 -7499
rect 65927 -7448 65979 -7438
rect 65786 -7490 65927 -7460
rect 65734 -7510 65786 -7500
rect 66118 -7448 66170 -7438
rect 65979 -7490 66118 -7460
rect 65927 -7510 65979 -7500
rect 66309 -7446 66361 -7436
rect 66170 -7490 66309 -7460
rect 66118 -7510 66170 -7500
rect 66504 -7448 66556 -7438
rect 66361 -7490 66504 -7460
rect 66309 -7508 66361 -7498
rect 66440 -7500 66504 -7490
rect 66440 -7510 66556 -7500
rect 66440 -7654 66510 -7510
rect 49940 -7664 66588 -7654
rect 47224 -7808 47652 -7752
rect 48274 -7706 48446 -7696
rect 48274 -7774 48446 -7764
rect 49940 -7766 66588 -7756
rect 68120 -7710 68292 -7700
rect 68120 -7778 68292 -7768
rect 68894 -7756 68924 -6672
rect 69290 -7756 69326 -6672
rect 68894 -7806 69326 -7756
rect 68584 -7808 69326 -7806
rect 47224 -8196 69326 -7808
rect 47482 -8198 69326 -8196
<< via2 >>
rect 48286 -5236 48444 -5178
rect 49920 -5280 66554 -5188
rect 68070 -5236 68228 -5178
rect 48274 -7764 48432 -7706
rect 49940 -7756 66574 -7664
rect 68120 -7768 68278 -7710
<< metal3 >>
rect 62104 -5160 62384 -5150
rect 67454 -5160 67734 -5150
rect 46340 -5178 69982 -5160
rect 46340 -5236 48286 -5178
rect 48444 -5188 68070 -5178
rect 48444 -5236 49920 -5188
rect 46340 -5280 49920 -5236
rect 66554 -5236 68070 -5188
rect 68228 -5236 69982 -5178
rect 66554 -5280 69982 -5236
rect 46340 -5438 69982 -5280
rect 49104 -6370 49384 -5438
rect 52114 -6370 52394 -5438
rect 55614 -6370 55894 -5438
rect 62104 -6370 62384 -5438
rect 64654 -6370 64934 -5438
rect 67454 -6370 67734 -5438
rect 46324 -6648 69966 -6370
rect 49104 -7510 49384 -6648
rect 52114 -7510 52394 -6648
rect 55614 -7510 55894 -6648
rect 62104 -7510 62384 -6648
rect 64654 -7510 64934 -6648
rect 67454 -7510 67734 -6648
rect 46350 -7664 69992 -7510
rect 46350 -7706 49940 -7664
rect 46350 -7764 48274 -7706
rect 48432 -7756 49940 -7706
rect 66574 -7710 69992 -7664
rect 66574 -7756 68120 -7710
rect 48432 -7764 68120 -7756
rect 46350 -7768 68120 -7764
rect 68278 -7768 69992 -7710
rect 46350 -7788 69992 -7768
use sky130_fd_pr__nfet_01v8_lvt_FKGFGD  XM20
timestamp 1662412052
transform 1 0 54905 0 1 -6780
box -3095 -310 3095 310
use sky130_fd_pr__nfet_01v8_lvt_FKGFGD  XM21
timestamp 1662412052
transform 1 0 54905 0 1 -6160
box -3095 -310 3095 310
use sky130_fd_pr__nfet_01v8_lvt_FKGFGD  XM22
timestamp 1662412052
transform 1 0 61095 0 1 -6160
box -3095 -310 3095 310
use sky130_fd_pr__nfet_01v8_lvt_FKGFGD  XM23
timestamp 1662412052
transform 1 0 61095 0 1 -6780
box -3095 -310 3095 310
use sky130_fd_pr__nfet_01v8_lvt_G3ZQK6  XM24
timestamp 1662412052
transform 1 0 58273 0 1 -5540
box -8423 -310 8423 310
use sky130_fd_pr__nfet_01v8_lvt_G3ZQK6  XM25
timestamp 1662412052
transform 1 0 58273 0 1 -7398
box -8423 -310 8423 310
use sky130_fd_pr__res_xhigh_po_5p73_4C7XCD  XR19
timestamp 1662952458
transform 0 1 47715 -1 0 -7211
box -739 -657 739 657
use sky130_fd_pr__res_xhigh_po_5p73_4C7XCD  XR20
timestamp 1662952458
transform 0 1 47715 -1 0 -5727
box -739 -657 739 657
use sky130_fd_pr__res_xhigh_po_5p73_QP6N54  XR21
timestamp 1662952458
transform 1 0 49111 0 1 -6518
box -739 -748 739 748
use sky130_fd_pr__res_xhigh_po_5p73_4C7XCD  XR22
timestamp 1662952458
transform 0 1 68837 -1 0 -5731
box -739 -657 739 657
use sky130_fd_pr__nfet_01v8_lvt_6H2JYD  sky130_fd_pr__nfet_01v8_lvt_6H2JYD_0
timestamp 1662976792
transform 0 1 51148 -1 0 -6469
box -211 -310 211 310
use sky130_fd_pr__nfet_01v8_lvt_6H2JYD  sky130_fd_pr__nfet_01v8_lvt_6H2JYD_1
timestamp 1662976792
transform 0 1 64558 -1 0 -6463
box -211 -310 211 310
use sky130_fd_pr__res_xhigh_po_5p73_4C7XCD  sky130_fd_pr__res_xhigh_po_5p73_4C7XCD_0
timestamp 1662952458
transform 0 1 68837 -1 0 -7211
box -739 -657 739 657
use sky130_fd_pr__res_xhigh_po_5p73_QP6N54  sky130_fd_pr__res_xhigh_po_5p73_QP6N54_0
timestamp 1662952458
transform 1 0 67439 0 1 -6468
box -739 -748 739 748
<< labels >>
rlabel metal3 46330 -6470 46330 -6470 7 vss
port 1 w
rlabel metal2 51160 -6220 51160 -6220 1 voutp
port 3 n
rlabel metal2 65180 -6220 65180 -6220 1 voutn
port 4 n
rlabel metal2 50660 -6720 50660 -6720 5 vd21
port 5 s
rlabel metal2 65770 -6710 65770 -6710 1 vd22
port 6 n
rlabel metal1 57930 -6930 57930 -6930 3 vinp
port 10 e
rlabel metal1 58070 -6930 58070 -6930 1 vinn
port 11 n
rlabel metal1 49890 -7550 49890 -7550 7 vc1
port 7 w
rlabel metal1 49880 -5390 49880 -5390 7 vc2
port 8 w
<< end >>
