magic
tech sky130A
magscale 1 2
timestamp 1671758665
<< nwell >>
rect -483 -4691 483 4691
<< pmoslvt >>
rect -287 2872 -187 4472
rect -129 2872 -29 4472
rect 29 2872 129 4472
rect 187 2872 287 4472
rect -287 1036 -187 2636
rect -129 1036 -29 2636
rect 29 1036 129 2636
rect 187 1036 287 2636
rect -287 -800 -187 800
rect -129 -800 -29 800
rect 29 -800 129 800
rect 187 -800 287 800
rect -287 -2636 -187 -1036
rect -129 -2636 -29 -1036
rect 29 -2636 129 -1036
rect 187 -2636 287 -1036
rect -287 -4472 -187 -2872
rect -129 -4472 -29 -2872
rect 29 -4472 129 -2872
rect 187 -4472 287 -2872
<< pdiff >>
rect -345 4460 -287 4472
rect -345 2884 -333 4460
rect -299 2884 -287 4460
rect -345 2872 -287 2884
rect -187 4460 -129 4472
rect -187 2884 -175 4460
rect -141 2884 -129 4460
rect -187 2872 -129 2884
rect -29 4460 29 4472
rect -29 2884 -17 4460
rect 17 2884 29 4460
rect -29 2872 29 2884
rect 129 4460 187 4472
rect 129 2884 141 4460
rect 175 2884 187 4460
rect 129 2872 187 2884
rect 287 4460 345 4472
rect 287 2884 299 4460
rect 333 2884 345 4460
rect 287 2872 345 2884
rect -345 2624 -287 2636
rect -345 1048 -333 2624
rect -299 1048 -287 2624
rect -345 1036 -287 1048
rect -187 2624 -129 2636
rect -187 1048 -175 2624
rect -141 1048 -129 2624
rect -187 1036 -129 1048
rect -29 2624 29 2636
rect -29 1048 -17 2624
rect 17 1048 29 2624
rect -29 1036 29 1048
rect 129 2624 187 2636
rect 129 1048 141 2624
rect 175 1048 187 2624
rect 129 1036 187 1048
rect 287 2624 345 2636
rect 287 1048 299 2624
rect 333 1048 345 2624
rect 287 1036 345 1048
rect -345 788 -287 800
rect -345 -788 -333 788
rect -299 -788 -287 788
rect -345 -800 -287 -788
rect -187 788 -129 800
rect -187 -788 -175 788
rect -141 -788 -129 788
rect -187 -800 -129 -788
rect -29 788 29 800
rect -29 -788 -17 788
rect 17 -788 29 788
rect -29 -800 29 -788
rect 129 788 187 800
rect 129 -788 141 788
rect 175 -788 187 788
rect 129 -800 187 -788
rect 287 788 345 800
rect 287 -788 299 788
rect 333 -788 345 788
rect 287 -800 345 -788
rect -345 -1048 -287 -1036
rect -345 -2624 -333 -1048
rect -299 -2624 -287 -1048
rect -345 -2636 -287 -2624
rect -187 -1048 -129 -1036
rect -187 -2624 -175 -1048
rect -141 -2624 -129 -1048
rect -187 -2636 -129 -2624
rect -29 -1048 29 -1036
rect -29 -2624 -17 -1048
rect 17 -2624 29 -1048
rect -29 -2636 29 -2624
rect 129 -1048 187 -1036
rect 129 -2624 141 -1048
rect 175 -2624 187 -1048
rect 129 -2636 187 -2624
rect 287 -1048 345 -1036
rect 287 -2624 299 -1048
rect 333 -2624 345 -1048
rect 287 -2636 345 -2624
rect -345 -2884 -287 -2872
rect -345 -4460 -333 -2884
rect -299 -4460 -287 -2884
rect -345 -4472 -287 -4460
rect -187 -2884 -129 -2872
rect -187 -4460 -175 -2884
rect -141 -4460 -129 -2884
rect -187 -4472 -129 -4460
rect -29 -2884 29 -2872
rect -29 -4460 -17 -2884
rect 17 -4460 29 -2884
rect -29 -4472 29 -4460
rect 129 -2884 187 -2872
rect 129 -4460 141 -2884
rect 175 -4460 187 -2884
rect 129 -4472 187 -4460
rect 287 -2884 345 -2872
rect 287 -4460 299 -2884
rect 333 -4460 345 -2884
rect 287 -4472 345 -4460
<< pdiffc >>
rect -333 2884 -299 4460
rect -175 2884 -141 4460
rect -17 2884 17 4460
rect 141 2884 175 4460
rect 299 2884 333 4460
rect -333 1048 -299 2624
rect -175 1048 -141 2624
rect -17 1048 17 2624
rect 141 1048 175 2624
rect 299 1048 333 2624
rect -333 -788 -299 788
rect -175 -788 -141 788
rect -17 -788 17 788
rect 141 -788 175 788
rect 299 -788 333 788
rect -333 -2624 -299 -1048
rect -175 -2624 -141 -1048
rect -17 -2624 17 -1048
rect 141 -2624 175 -1048
rect 299 -2624 333 -1048
rect -333 -4460 -299 -2884
rect -175 -4460 -141 -2884
rect -17 -4460 17 -2884
rect 141 -4460 175 -2884
rect 299 -4460 333 -2884
<< nsubdiff >>
rect -447 4621 -351 4655
rect 351 4621 447 4655
rect -447 -4621 -413 4621
rect 413 -4621 447 4621
rect -447 -4655 -351 -4621
rect 351 -4655 447 -4621
<< nsubdiffcont >>
rect -351 4621 351 4655
rect -351 -4655 351 -4621
<< poly >>
rect -287 4553 -187 4569
rect -287 4519 -271 4553
rect -203 4519 -187 4553
rect -287 4472 -187 4519
rect -129 4553 -29 4569
rect -129 4519 -113 4553
rect -45 4519 -29 4553
rect -129 4472 -29 4519
rect 29 4553 129 4569
rect 29 4519 45 4553
rect 113 4519 129 4553
rect 29 4472 129 4519
rect 187 4553 287 4569
rect 187 4519 203 4553
rect 271 4519 287 4553
rect 187 4472 287 4519
rect -287 2825 -187 2872
rect -287 2791 -271 2825
rect -203 2791 -187 2825
rect -287 2775 -187 2791
rect -129 2825 -29 2872
rect -129 2791 -113 2825
rect -45 2791 -29 2825
rect -129 2775 -29 2791
rect 29 2825 129 2872
rect 29 2791 45 2825
rect 113 2791 129 2825
rect 29 2775 129 2791
rect 187 2825 287 2872
rect 187 2791 203 2825
rect 271 2791 287 2825
rect 187 2775 287 2791
rect -287 2717 -187 2733
rect -287 2683 -271 2717
rect -203 2683 -187 2717
rect -287 2636 -187 2683
rect -129 2717 -29 2733
rect -129 2683 -113 2717
rect -45 2683 -29 2717
rect -129 2636 -29 2683
rect 29 2717 129 2733
rect 29 2683 45 2717
rect 113 2683 129 2717
rect 29 2636 129 2683
rect 187 2717 287 2733
rect 187 2683 203 2717
rect 271 2683 287 2717
rect 187 2636 287 2683
rect -287 989 -187 1036
rect -287 955 -271 989
rect -203 955 -187 989
rect -287 939 -187 955
rect -129 989 -29 1036
rect -129 955 -113 989
rect -45 955 -29 989
rect -129 939 -29 955
rect 29 989 129 1036
rect 29 955 45 989
rect 113 955 129 989
rect 29 939 129 955
rect 187 989 287 1036
rect 187 955 203 989
rect 271 955 287 989
rect 187 939 287 955
rect -287 881 -187 897
rect -287 847 -271 881
rect -203 847 -187 881
rect -287 800 -187 847
rect -129 881 -29 897
rect -129 847 -113 881
rect -45 847 -29 881
rect -129 800 -29 847
rect 29 881 129 897
rect 29 847 45 881
rect 113 847 129 881
rect 29 800 129 847
rect 187 881 287 897
rect 187 847 203 881
rect 271 847 287 881
rect 187 800 287 847
rect -287 -847 -187 -800
rect -287 -881 -271 -847
rect -203 -881 -187 -847
rect -287 -897 -187 -881
rect -129 -847 -29 -800
rect -129 -881 -113 -847
rect -45 -881 -29 -847
rect -129 -897 -29 -881
rect 29 -847 129 -800
rect 29 -881 45 -847
rect 113 -881 129 -847
rect 29 -897 129 -881
rect 187 -847 287 -800
rect 187 -881 203 -847
rect 271 -881 287 -847
rect 187 -897 287 -881
rect -287 -955 -187 -939
rect -287 -989 -271 -955
rect -203 -989 -187 -955
rect -287 -1036 -187 -989
rect -129 -955 -29 -939
rect -129 -989 -113 -955
rect -45 -989 -29 -955
rect -129 -1036 -29 -989
rect 29 -955 129 -939
rect 29 -989 45 -955
rect 113 -989 129 -955
rect 29 -1036 129 -989
rect 187 -955 287 -939
rect 187 -989 203 -955
rect 271 -989 287 -955
rect 187 -1036 287 -989
rect -287 -2683 -187 -2636
rect -287 -2717 -271 -2683
rect -203 -2717 -187 -2683
rect -287 -2733 -187 -2717
rect -129 -2683 -29 -2636
rect -129 -2717 -113 -2683
rect -45 -2717 -29 -2683
rect -129 -2733 -29 -2717
rect 29 -2683 129 -2636
rect 29 -2717 45 -2683
rect 113 -2717 129 -2683
rect 29 -2733 129 -2717
rect 187 -2683 287 -2636
rect 187 -2717 203 -2683
rect 271 -2717 287 -2683
rect 187 -2733 287 -2717
rect -287 -2791 -187 -2775
rect -287 -2825 -271 -2791
rect -203 -2825 -187 -2791
rect -287 -2872 -187 -2825
rect -129 -2791 -29 -2775
rect -129 -2825 -113 -2791
rect -45 -2825 -29 -2791
rect -129 -2872 -29 -2825
rect 29 -2791 129 -2775
rect 29 -2825 45 -2791
rect 113 -2825 129 -2791
rect 29 -2872 129 -2825
rect 187 -2791 287 -2775
rect 187 -2825 203 -2791
rect 271 -2825 287 -2791
rect 187 -2872 287 -2825
rect -287 -4519 -187 -4472
rect -287 -4553 -271 -4519
rect -203 -4553 -187 -4519
rect -287 -4569 -187 -4553
rect -129 -4519 -29 -4472
rect -129 -4553 -113 -4519
rect -45 -4553 -29 -4519
rect -129 -4569 -29 -4553
rect 29 -4519 129 -4472
rect 29 -4553 45 -4519
rect 113 -4553 129 -4519
rect 29 -4569 129 -4553
rect 187 -4519 287 -4472
rect 187 -4553 203 -4519
rect 271 -4553 287 -4519
rect 187 -4569 287 -4553
<< polycont >>
rect -271 4519 -203 4553
rect -113 4519 -45 4553
rect 45 4519 113 4553
rect 203 4519 271 4553
rect -271 2791 -203 2825
rect -113 2791 -45 2825
rect 45 2791 113 2825
rect 203 2791 271 2825
rect -271 2683 -203 2717
rect -113 2683 -45 2717
rect 45 2683 113 2717
rect 203 2683 271 2717
rect -271 955 -203 989
rect -113 955 -45 989
rect 45 955 113 989
rect 203 955 271 989
rect -271 847 -203 881
rect -113 847 -45 881
rect 45 847 113 881
rect 203 847 271 881
rect -271 -881 -203 -847
rect -113 -881 -45 -847
rect 45 -881 113 -847
rect 203 -881 271 -847
rect -271 -989 -203 -955
rect -113 -989 -45 -955
rect 45 -989 113 -955
rect 203 -989 271 -955
rect -271 -2717 -203 -2683
rect -113 -2717 -45 -2683
rect 45 -2717 113 -2683
rect 203 -2717 271 -2683
rect -271 -2825 -203 -2791
rect -113 -2825 -45 -2791
rect 45 -2825 113 -2791
rect 203 -2825 271 -2791
rect -271 -4553 -203 -4519
rect -113 -4553 -45 -4519
rect 45 -4553 113 -4519
rect 203 -4553 271 -4519
<< locali >>
rect -447 4621 -351 4655
rect 351 4621 447 4655
rect -447 -4621 -413 4621
rect -287 4519 -271 4553
rect -203 4519 -187 4553
rect -129 4519 -113 4553
rect -45 4519 -29 4553
rect 29 4519 45 4553
rect 113 4519 129 4553
rect 187 4519 203 4553
rect 271 4519 287 4553
rect -333 4460 -299 4476
rect -333 2868 -299 2884
rect -175 4460 -141 4476
rect -175 2868 -141 2884
rect -17 4460 17 4476
rect -17 2868 17 2884
rect 141 4460 175 4476
rect 141 2868 175 2884
rect 299 4460 333 4476
rect 299 2868 333 2884
rect -287 2791 -271 2825
rect -203 2791 -187 2825
rect -129 2791 -113 2825
rect -45 2791 -29 2825
rect 29 2791 45 2825
rect 113 2791 129 2825
rect 187 2791 203 2825
rect 271 2791 287 2825
rect -287 2683 -271 2717
rect -203 2683 -187 2717
rect -129 2683 -113 2717
rect -45 2683 -29 2717
rect 29 2683 45 2717
rect 113 2683 129 2717
rect 187 2683 203 2717
rect 271 2683 287 2717
rect -333 2624 -299 2640
rect -333 1032 -299 1048
rect -175 2624 -141 2640
rect -175 1032 -141 1048
rect -17 2624 17 2640
rect -17 1032 17 1048
rect 141 2624 175 2640
rect 141 1032 175 1048
rect 299 2624 333 2640
rect 299 1032 333 1048
rect -287 955 -271 989
rect -203 955 -187 989
rect -129 955 -113 989
rect -45 955 -29 989
rect 29 955 45 989
rect 113 955 129 989
rect 187 955 203 989
rect 271 955 287 989
rect -287 847 -271 881
rect -203 847 -187 881
rect -129 847 -113 881
rect -45 847 -29 881
rect 29 847 45 881
rect 113 847 129 881
rect 187 847 203 881
rect 271 847 287 881
rect -333 788 -299 804
rect -333 -804 -299 -788
rect -175 788 -141 804
rect -175 -804 -141 -788
rect -17 788 17 804
rect -17 -804 17 -788
rect 141 788 175 804
rect 141 -804 175 -788
rect 299 788 333 804
rect 299 -804 333 -788
rect -287 -881 -271 -847
rect -203 -881 -187 -847
rect -129 -881 -113 -847
rect -45 -881 -29 -847
rect 29 -881 45 -847
rect 113 -881 129 -847
rect 187 -881 203 -847
rect 271 -881 287 -847
rect -287 -989 -271 -955
rect -203 -989 -187 -955
rect -129 -989 -113 -955
rect -45 -989 -29 -955
rect 29 -989 45 -955
rect 113 -989 129 -955
rect 187 -989 203 -955
rect 271 -989 287 -955
rect -333 -1048 -299 -1032
rect -333 -2640 -299 -2624
rect -175 -1048 -141 -1032
rect -175 -2640 -141 -2624
rect -17 -1048 17 -1032
rect -17 -2640 17 -2624
rect 141 -1048 175 -1032
rect 141 -2640 175 -2624
rect 299 -1048 333 -1032
rect 299 -2640 333 -2624
rect -287 -2717 -271 -2683
rect -203 -2717 -187 -2683
rect -129 -2717 -113 -2683
rect -45 -2717 -29 -2683
rect 29 -2717 45 -2683
rect 113 -2717 129 -2683
rect 187 -2717 203 -2683
rect 271 -2717 287 -2683
rect -287 -2825 -271 -2791
rect -203 -2825 -187 -2791
rect -129 -2825 -113 -2791
rect -45 -2825 -29 -2791
rect 29 -2825 45 -2791
rect 113 -2825 129 -2791
rect 187 -2825 203 -2791
rect 271 -2825 287 -2791
rect -333 -2884 -299 -2868
rect -333 -4476 -299 -4460
rect -175 -2884 -141 -2868
rect -175 -4476 -141 -4460
rect -17 -2884 17 -2868
rect -17 -4476 17 -4460
rect 141 -2884 175 -2868
rect 141 -4476 175 -4460
rect 299 -2884 333 -2868
rect 299 -4476 333 -4460
rect -287 -4553 -271 -4519
rect -203 -4553 -187 -4519
rect -129 -4553 -113 -4519
rect -45 -4553 -29 -4519
rect 29 -4553 45 -4519
rect 113 -4553 129 -4519
rect 187 -4553 203 -4519
rect 271 -4553 287 -4519
rect 413 -4621 447 4621
rect -447 -4655 -351 -4621
rect 351 -4655 447 -4621
<< viali >>
rect -271 4519 -203 4553
rect -113 4519 -45 4553
rect 45 4519 113 4553
rect 203 4519 271 4553
rect -333 2884 -299 4460
rect -175 2884 -141 4460
rect -17 2884 17 4460
rect 141 2884 175 4460
rect 299 2884 333 4460
rect -271 2791 -203 2825
rect -113 2791 -45 2825
rect 45 2791 113 2825
rect 203 2791 271 2825
rect -271 2683 -203 2717
rect -113 2683 -45 2717
rect 45 2683 113 2717
rect 203 2683 271 2717
rect -333 1048 -299 2624
rect -175 1048 -141 2624
rect -17 1048 17 2624
rect 141 1048 175 2624
rect 299 1048 333 2624
rect -271 955 -203 989
rect -113 955 -45 989
rect 45 955 113 989
rect 203 955 271 989
rect -271 847 -203 881
rect -113 847 -45 881
rect 45 847 113 881
rect 203 847 271 881
rect -333 -788 -299 788
rect -175 -788 -141 788
rect -17 -788 17 788
rect 141 -788 175 788
rect 299 -788 333 788
rect -271 -881 -203 -847
rect -113 -881 -45 -847
rect 45 -881 113 -847
rect 203 -881 271 -847
rect -271 -989 -203 -955
rect -113 -989 -45 -955
rect 45 -989 113 -955
rect 203 -989 271 -955
rect -333 -2624 -299 -1048
rect -175 -2624 -141 -1048
rect -17 -2624 17 -1048
rect 141 -2624 175 -1048
rect 299 -2624 333 -1048
rect -271 -2717 -203 -2683
rect -113 -2717 -45 -2683
rect 45 -2717 113 -2683
rect 203 -2717 271 -2683
rect -271 -2825 -203 -2791
rect -113 -2825 -45 -2791
rect 45 -2825 113 -2791
rect 203 -2825 271 -2791
rect -333 -4460 -299 -2884
rect -175 -4460 -141 -2884
rect -17 -4460 17 -2884
rect 141 -4460 175 -2884
rect 299 -4460 333 -2884
rect -271 -4553 -203 -4519
rect -113 -4553 -45 -4519
rect 45 -4553 113 -4519
rect 203 -4553 271 -4519
<< metal1 >>
rect -283 4553 -191 4559
rect -283 4519 -271 4553
rect -203 4519 -191 4553
rect -283 4513 -191 4519
rect -125 4553 -33 4559
rect -125 4519 -113 4553
rect -45 4519 -33 4553
rect -125 4513 -33 4519
rect 33 4553 125 4559
rect 33 4519 45 4553
rect 113 4519 125 4553
rect 33 4513 125 4519
rect 191 4553 283 4559
rect 191 4519 203 4553
rect 271 4519 283 4553
rect 191 4513 283 4519
rect -339 4460 -293 4472
rect -339 2884 -333 4460
rect -299 2884 -293 4460
rect -339 2872 -293 2884
rect -181 4460 -135 4472
rect -181 2884 -175 4460
rect -141 2884 -135 4460
rect -181 2872 -135 2884
rect -23 4460 23 4472
rect -23 2884 -17 4460
rect 17 2884 23 4460
rect -23 2872 23 2884
rect 135 4460 181 4472
rect 135 2884 141 4460
rect 175 2884 181 4460
rect 135 2872 181 2884
rect 293 4460 339 4472
rect 293 2884 299 4460
rect 333 2884 339 4460
rect 293 2872 339 2884
rect -283 2825 -191 2831
rect -283 2791 -271 2825
rect -203 2791 -191 2825
rect -283 2785 -191 2791
rect -125 2825 -33 2831
rect -125 2791 -113 2825
rect -45 2791 -33 2825
rect -125 2785 -33 2791
rect 33 2825 125 2831
rect 33 2791 45 2825
rect 113 2791 125 2825
rect 33 2785 125 2791
rect 191 2825 283 2831
rect 191 2791 203 2825
rect 271 2791 283 2825
rect 191 2785 283 2791
rect -283 2717 -191 2723
rect -283 2683 -271 2717
rect -203 2683 -191 2717
rect -283 2677 -191 2683
rect -125 2717 -33 2723
rect -125 2683 -113 2717
rect -45 2683 -33 2717
rect -125 2677 -33 2683
rect 33 2717 125 2723
rect 33 2683 45 2717
rect 113 2683 125 2717
rect 33 2677 125 2683
rect 191 2717 283 2723
rect 191 2683 203 2717
rect 271 2683 283 2717
rect 191 2677 283 2683
rect -339 2624 -293 2636
rect -339 1048 -333 2624
rect -299 1048 -293 2624
rect -339 1036 -293 1048
rect -181 2624 -135 2636
rect -181 1048 -175 2624
rect -141 1048 -135 2624
rect -181 1036 -135 1048
rect -23 2624 23 2636
rect -23 1048 -17 2624
rect 17 1048 23 2624
rect -23 1036 23 1048
rect 135 2624 181 2636
rect 135 1048 141 2624
rect 175 1048 181 2624
rect 135 1036 181 1048
rect 293 2624 339 2636
rect 293 1048 299 2624
rect 333 1048 339 2624
rect 293 1036 339 1048
rect -283 989 -191 995
rect -283 955 -271 989
rect -203 955 -191 989
rect -283 949 -191 955
rect -125 989 -33 995
rect -125 955 -113 989
rect -45 955 -33 989
rect -125 949 -33 955
rect 33 989 125 995
rect 33 955 45 989
rect 113 955 125 989
rect 33 949 125 955
rect 191 989 283 995
rect 191 955 203 989
rect 271 955 283 989
rect 191 949 283 955
rect -283 881 -191 887
rect -283 847 -271 881
rect -203 847 -191 881
rect -283 841 -191 847
rect -125 881 -33 887
rect -125 847 -113 881
rect -45 847 -33 881
rect -125 841 -33 847
rect 33 881 125 887
rect 33 847 45 881
rect 113 847 125 881
rect 33 841 125 847
rect 191 881 283 887
rect 191 847 203 881
rect 271 847 283 881
rect 191 841 283 847
rect -339 788 -293 800
rect -339 -788 -333 788
rect -299 -788 -293 788
rect -339 -800 -293 -788
rect -181 788 -135 800
rect -181 -788 -175 788
rect -141 -788 -135 788
rect -181 -800 -135 -788
rect -23 788 23 800
rect -23 -788 -17 788
rect 17 -788 23 788
rect -23 -800 23 -788
rect 135 788 181 800
rect 135 -788 141 788
rect 175 -788 181 788
rect 135 -800 181 -788
rect 293 788 339 800
rect 293 -788 299 788
rect 333 -788 339 788
rect 293 -800 339 -788
rect -283 -847 -191 -841
rect -283 -881 -271 -847
rect -203 -881 -191 -847
rect -283 -887 -191 -881
rect -125 -847 -33 -841
rect -125 -881 -113 -847
rect -45 -881 -33 -847
rect -125 -887 -33 -881
rect 33 -847 125 -841
rect 33 -881 45 -847
rect 113 -881 125 -847
rect 33 -887 125 -881
rect 191 -847 283 -841
rect 191 -881 203 -847
rect 271 -881 283 -847
rect 191 -887 283 -881
rect -283 -955 -191 -949
rect -283 -989 -271 -955
rect -203 -989 -191 -955
rect -283 -995 -191 -989
rect -125 -955 -33 -949
rect -125 -989 -113 -955
rect -45 -989 -33 -955
rect -125 -995 -33 -989
rect 33 -955 125 -949
rect 33 -989 45 -955
rect 113 -989 125 -955
rect 33 -995 125 -989
rect 191 -955 283 -949
rect 191 -989 203 -955
rect 271 -989 283 -955
rect 191 -995 283 -989
rect -339 -1048 -293 -1036
rect -339 -2624 -333 -1048
rect -299 -2624 -293 -1048
rect -339 -2636 -293 -2624
rect -181 -1048 -135 -1036
rect -181 -2624 -175 -1048
rect -141 -2624 -135 -1048
rect -181 -2636 -135 -2624
rect -23 -1048 23 -1036
rect -23 -2624 -17 -1048
rect 17 -2624 23 -1048
rect -23 -2636 23 -2624
rect 135 -1048 181 -1036
rect 135 -2624 141 -1048
rect 175 -2624 181 -1048
rect 135 -2636 181 -2624
rect 293 -1048 339 -1036
rect 293 -2624 299 -1048
rect 333 -2624 339 -1048
rect 293 -2636 339 -2624
rect -283 -2683 -191 -2677
rect -283 -2717 -271 -2683
rect -203 -2717 -191 -2683
rect -283 -2723 -191 -2717
rect -125 -2683 -33 -2677
rect -125 -2717 -113 -2683
rect -45 -2717 -33 -2683
rect -125 -2723 -33 -2717
rect 33 -2683 125 -2677
rect 33 -2717 45 -2683
rect 113 -2717 125 -2683
rect 33 -2723 125 -2717
rect 191 -2683 283 -2677
rect 191 -2717 203 -2683
rect 271 -2717 283 -2683
rect 191 -2723 283 -2717
rect -283 -2791 -191 -2785
rect -283 -2825 -271 -2791
rect -203 -2825 -191 -2791
rect -283 -2831 -191 -2825
rect -125 -2791 -33 -2785
rect -125 -2825 -113 -2791
rect -45 -2825 -33 -2791
rect -125 -2831 -33 -2825
rect 33 -2791 125 -2785
rect 33 -2825 45 -2791
rect 113 -2825 125 -2791
rect 33 -2831 125 -2825
rect 191 -2791 283 -2785
rect 191 -2825 203 -2791
rect 271 -2825 283 -2791
rect 191 -2831 283 -2825
rect -339 -2884 -293 -2872
rect -339 -4460 -333 -2884
rect -299 -4460 -293 -2884
rect -339 -4472 -293 -4460
rect -181 -2884 -135 -2872
rect -181 -4460 -175 -2884
rect -141 -4460 -135 -2884
rect -181 -4472 -135 -4460
rect -23 -2884 23 -2872
rect -23 -4460 -17 -2884
rect 17 -4460 23 -2884
rect -23 -4472 23 -4460
rect 135 -2884 181 -2872
rect 135 -4460 141 -2884
rect 175 -4460 181 -2884
rect 135 -4472 181 -4460
rect 293 -2884 339 -2872
rect 293 -4460 299 -2884
rect 333 -4460 339 -2884
rect 293 -4472 339 -4460
rect -283 -4519 -191 -4513
rect -283 -4553 -271 -4519
rect -203 -4553 -191 -4519
rect -283 -4559 -191 -4553
rect -125 -4519 -33 -4513
rect -125 -4553 -113 -4519
rect -45 -4553 -33 -4519
rect -125 -4559 -33 -4553
rect 33 -4519 125 -4513
rect 33 -4553 45 -4519
rect 113 -4553 125 -4519
rect 33 -4559 125 -4553
rect 191 -4519 283 -4513
rect 191 -4553 203 -4519
rect 271 -4553 283 -4519
rect 191 -4559 283 -4553
<< properties >>
string FIXED_BBOX -430 -4638 430 4638
string gencell sky130_fd_pr__pfet_01v8_lvt
string library sky130
string parameters w 8 l 0.5 m 5 nf 4 diffcov 100 polycov 100 guard 1 glc 0 grc 0 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.35 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
