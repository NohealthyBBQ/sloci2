magic
tech sky130A
magscale 1 2
timestamp 1660068957
<< error_p >>
rect -2847 181 -2785 187
rect -2719 181 -2657 187
rect -2591 181 -2529 187
rect -2463 181 -2401 187
rect -2335 181 -2273 187
rect -2207 181 -2145 187
rect -2079 181 -2017 187
rect -1951 181 -1889 187
rect -1823 181 -1761 187
rect -1695 181 -1633 187
rect -1567 181 -1505 187
rect -1439 181 -1377 187
rect -1311 181 -1249 187
rect -1183 181 -1121 187
rect -1055 181 -993 187
rect -927 181 -865 187
rect -799 181 -737 187
rect -671 181 -609 187
rect -543 181 -481 187
rect -415 181 -353 187
rect -287 181 -225 187
rect -159 181 -97 187
rect -31 181 31 187
rect 97 181 159 187
rect 225 181 287 187
rect 353 181 415 187
rect 481 181 543 187
rect 609 181 671 187
rect 737 181 799 187
rect 865 181 927 187
rect 993 181 1055 187
rect 1121 181 1183 187
rect 1249 181 1311 187
rect 1377 181 1439 187
rect 1505 181 1567 187
rect 1633 181 1695 187
rect 1761 181 1823 187
rect 1889 181 1951 187
rect 2017 181 2079 187
rect 2145 181 2207 187
rect 2273 181 2335 187
rect 2401 181 2463 187
rect 2529 181 2591 187
rect 2657 181 2719 187
rect 2785 181 2847 187
rect -2847 147 -2835 181
rect -2719 147 -2707 181
rect -2591 147 -2579 181
rect -2463 147 -2451 181
rect -2335 147 -2323 181
rect -2207 147 -2195 181
rect -2079 147 -2067 181
rect -1951 147 -1939 181
rect -1823 147 -1811 181
rect -1695 147 -1683 181
rect -1567 147 -1555 181
rect -1439 147 -1427 181
rect -1311 147 -1299 181
rect -1183 147 -1171 181
rect -1055 147 -1043 181
rect -927 147 -915 181
rect -799 147 -787 181
rect -671 147 -659 181
rect -543 147 -531 181
rect -415 147 -403 181
rect -287 147 -275 181
rect -159 147 -147 181
rect -31 147 -19 181
rect 97 147 109 181
rect 225 147 237 181
rect 353 147 365 181
rect 481 147 493 181
rect 609 147 621 181
rect 737 147 749 181
rect 865 147 877 181
rect 993 147 1005 181
rect 1121 147 1133 181
rect 1249 147 1261 181
rect 1377 147 1389 181
rect 1505 147 1517 181
rect 1633 147 1645 181
rect 1761 147 1773 181
rect 1889 147 1901 181
rect 2017 147 2029 181
rect 2145 147 2157 181
rect 2273 147 2285 181
rect 2401 147 2413 181
rect 2529 147 2541 181
rect 2657 147 2669 181
rect 2785 147 2797 181
rect -2847 141 -2785 147
rect -2719 141 -2657 147
rect -2591 141 -2529 147
rect -2463 141 -2401 147
rect -2335 141 -2273 147
rect -2207 141 -2145 147
rect -2079 141 -2017 147
rect -1951 141 -1889 147
rect -1823 141 -1761 147
rect -1695 141 -1633 147
rect -1567 141 -1505 147
rect -1439 141 -1377 147
rect -1311 141 -1249 147
rect -1183 141 -1121 147
rect -1055 141 -993 147
rect -927 141 -865 147
rect -799 141 -737 147
rect -671 141 -609 147
rect -543 141 -481 147
rect -415 141 -353 147
rect -287 141 -225 147
rect -159 141 -97 147
rect -31 141 31 147
rect 97 141 159 147
rect 225 141 287 147
rect 353 141 415 147
rect 481 141 543 147
rect 609 141 671 147
rect 737 141 799 147
rect 865 141 927 147
rect 993 141 1055 147
rect 1121 141 1183 147
rect 1249 141 1311 147
rect 1377 141 1439 147
rect 1505 141 1567 147
rect 1633 141 1695 147
rect 1761 141 1823 147
rect 1889 141 1951 147
rect 2017 141 2079 147
rect 2145 141 2207 147
rect 2273 141 2335 147
rect 2401 141 2463 147
rect 2529 141 2591 147
rect 2657 141 2719 147
rect 2785 141 2847 147
rect -2847 -147 -2785 -141
rect -2719 -147 -2657 -141
rect -2591 -147 -2529 -141
rect -2463 -147 -2401 -141
rect -2335 -147 -2273 -141
rect -2207 -147 -2145 -141
rect -2079 -147 -2017 -141
rect -1951 -147 -1889 -141
rect -1823 -147 -1761 -141
rect -1695 -147 -1633 -141
rect -1567 -147 -1505 -141
rect -1439 -147 -1377 -141
rect -1311 -147 -1249 -141
rect -1183 -147 -1121 -141
rect -1055 -147 -993 -141
rect -927 -147 -865 -141
rect -799 -147 -737 -141
rect -671 -147 -609 -141
rect -543 -147 -481 -141
rect -415 -147 -353 -141
rect -287 -147 -225 -141
rect -159 -147 -97 -141
rect -31 -147 31 -141
rect 97 -147 159 -141
rect 225 -147 287 -141
rect 353 -147 415 -141
rect 481 -147 543 -141
rect 609 -147 671 -141
rect 737 -147 799 -141
rect 865 -147 927 -141
rect 993 -147 1055 -141
rect 1121 -147 1183 -141
rect 1249 -147 1311 -141
rect 1377 -147 1439 -141
rect 1505 -147 1567 -141
rect 1633 -147 1695 -141
rect 1761 -147 1823 -141
rect 1889 -147 1951 -141
rect 2017 -147 2079 -141
rect 2145 -147 2207 -141
rect 2273 -147 2335 -141
rect 2401 -147 2463 -141
rect 2529 -147 2591 -141
rect 2657 -147 2719 -141
rect 2785 -147 2847 -141
rect -2847 -181 -2835 -147
rect -2719 -181 -2707 -147
rect -2591 -181 -2579 -147
rect -2463 -181 -2451 -147
rect -2335 -181 -2323 -147
rect -2207 -181 -2195 -147
rect -2079 -181 -2067 -147
rect -1951 -181 -1939 -147
rect -1823 -181 -1811 -147
rect -1695 -181 -1683 -147
rect -1567 -181 -1555 -147
rect -1439 -181 -1427 -147
rect -1311 -181 -1299 -147
rect -1183 -181 -1171 -147
rect -1055 -181 -1043 -147
rect -927 -181 -915 -147
rect -799 -181 -787 -147
rect -671 -181 -659 -147
rect -543 -181 -531 -147
rect -415 -181 -403 -147
rect -287 -181 -275 -147
rect -159 -181 -147 -147
rect -31 -181 -19 -147
rect 97 -181 109 -147
rect 225 -181 237 -147
rect 353 -181 365 -147
rect 481 -181 493 -147
rect 609 -181 621 -147
rect 737 -181 749 -147
rect 865 -181 877 -147
rect 993 -181 1005 -147
rect 1121 -181 1133 -147
rect 1249 -181 1261 -147
rect 1377 -181 1389 -147
rect 1505 -181 1517 -147
rect 1633 -181 1645 -147
rect 1761 -181 1773 -147
rect 1889 -181 1901 -147
rect 2017 -181 2029 -147
rect 2145 -181 2157 -147
rect 2273 -181 2285 -147
rect 2401 -181 2413 -147
rect 2529 -181 2541 -147
rect 2657 -181 2669 -147
rect 2785 -181 2797 -147
rect -2847 -187 -2785 -181
rect -2719 -187 -2657 -181
rect -2591 -187 -2529 -181
rect -2463 -187 -2401 -181
rect -2335 -187 -2273 -181
rect -2207 -187 -2145 -181
rect -2079 -187 -2017 -181
rect -1951 -187 -1889 -181
rect -1823 -187 -1761 -181
rect -1695 -187 -1633 -181
rect -1567 -187 -1505 -181
rect -1439 -187 -1377 -181
rect -1311 -187 -1249 -181
rect -1183 -187 -1121 -181
rect -1055 -187 -993 -181
rect -927 -187 -865 -181
rect -799 -187 -737 -181
rect -671 -187 -609 -181
rect -543 -187 -481 -181
rect -415 -187 -353 -181
rect -287 -187 -225 -181
rect -159 -187 -97 -181
rect -31 -187 31 -181
rect 97 -187 159 -181
rect 225 -187 287 -181
rect 353 -187 415 -181
rect 481 -187 543 -181
rect 609 -187 671 -181
rect 737 -187 799 -181
rect 865 -187 927 -181
rect 993 -187 1055 -181
rect 1121 -187 1183 -181
rect 1249 -187 1311 -181
rect 1377 -187 1439 -181
rect 1505 -187 1567 -181
rect 1633 -187 1695 -181
rect 1761 -187 1823 -181
rect 1889 -187 1951 -181
rect 2017 -187 2079 -181
rect 2145 -187 2207 -181
rect 2273 -187 2335 -181
rect 2401 -187 2463 -181
rect 2529 -187 2591 -181
rect 2657 -187 2719 -181
rect 2785 -187 2847 -181
<< nwell >>
rect -3047 -319 3047 319
<< pmoslvt >>
rect -2851 -100 -2781 100
rect -2723 -100 -2653 100
rect -2595 -100 -2525 100
rect -2467 -100 -2397 100
rect -2339 -100 -2269 100
rect -2211 -100 -2141 100
rect -2083 -100 -2013 100
rect -1955 -100 -1885 100
rect -1827 -100 -1757 100
rect -1699 -100 -1629 100
rect -1571 -100 -1501 100
rect -1443 -100 -1373 100
rect -1315 -100 -1245 100
rect -1187 -100 -1117 100
rect -1059 -100 -989 100
rect -931 -100 -861 100
rect -803 -100 -733 100
rect -675 -100 -605 100
rect -547 -100 -477 100
rect -419 -100 -349 100
rect -291 -100 -221 100
rect -163 -100 -93 100
rect -35 -100 35 100
rect 93 -100 163 100
rect 221 -100 291 100
rect 349 -100 419 100
rect 477 -100 547 100
rect 605 -100 675 100
rect 733 -100 803 100
rect 861 -100 931 100
rect 989 -100 1059 100
rect 1117 -100 1187 100
rect 1245 -100 1315 100
rect 1373 -100 1443 100
rect 1501 -100 1571 100
rect 1629 -100 1699 100
rect 1757 -100 1827 100
rect 1885 -100 1955 100
rect 2013 -100 2083 100
rect 2141 -100 2211 100
rect 2269 -100 2339 100
rect 2397 -100 2467 100
rect 2525 -100 2595 100
rect 2653 -100 2723 100
rect 2781 -100 2851 100
<< pdiff >>
rect -2909 88 -2851 100
rect -2909 -88 -2897 88
rect -2863 -88 -2851 88
rect -2909 -100 -2851 -88
rect -2781 88 -2723 100
rect -2781 -88 -2769 88
rect -2735 -88 -2723 88
rect -2781 -100 -2723 -88
rect -2653 88 -2595 100
rect -2653 -88 -2641 88
rect -2607 -88 -2595 88
rect -2653 -100 -2595 -88
rect -2525 88 -2467 100
rect -2525 -88 -2513 88
rect -2479 -88 -2467 88
rect -2525 -100 -2467 -88
rect -2397 88 -2339 100
rect -2397 -88 -2385 88
rect -2351 -88 -2339 88
rect -2397 -100 -2339 -88
rect -2269 88 -2211 100
rect -2269 -88 -2257 88
rect -2223 -88 -2211 88
rect -2269 -100 -2211 -88
rect -2141 88 -2083 100
rect -2141 -88 -2129 88
rect -2095 -88 -2083 88
rect -2141 -100 -2083 -88
rect -2013 88 -1955 100
rect -2013 -88 -2001 88
rect -1967 -88 -1955 88
rect -2013 -100 -1955 -88
rect -1885 88 -1827 100
rect -1885 -88 -1873 88
rect -1839 -88 -1827 88
rect -1885 -100 -1827 -88
rect -1757 88 -1699 100
rect -1757 -88 -1745 88
rect -1711 -88 -1699 88
rect -1757 -100 -1699 -88
rect -1629 88 -1571 100
rect -1629 -88 -1617 88
rect -1583 -88 -1571 88
rect -1629 -100 -1571 -88
rect -1501 88 -1443 100
rect -1501 -88 -1489 88
rect -1455 -88 -1443 88
rect -1501 -100 -1443 -88
rect -1373 88 -1315 100
rect -1373 -88 -1361 88
rect -1327 -88 -1315 88
rect -1373 -100 -1315 -88
rect -1245 88 -1187 100
rect -1245 -88 -1233 88
rect -1199 -88 -1187 88
rect -1245 -100 -1187 -88
rect -1117 88 -1059 100
rect -1117 -88 -1105 88
rect -1071 -88 -1059 88
rect -1117 -100 -1059 -88
rect -989 88 -931 100
rect -989 -88 -977 88
rect -943 -88 -931 88
rect -989 -100 -931 -88
rect -861 88 -803 100
rect -861 -88 -849 88
rect -815 -88 -803 88
rect -861 -100 -803 -88
rect -733 88 -675 100
rect -733 -88 -721 88
rect -687 -88 -675 88
rect -733 -100 -675 -88
rect -605 88 -547 100
rect -605 -88 -593 88
rect -559 -88 -547 88
rect -605 -100 -547 -88
rect -477 88 -419 100
rect -477 -88 -465 88
rect -431 -88 -419 88
rect -477 -100 -419 -88
rect -349 88 -291 100
rect -349 -88 -337 88
rect -303 -88 -291 88
rect -349 -100 -291 -88
rect -221 88 -163 100
rect -221 -88 -209 88
rect -175 -88 -163 88
rect -221 -100 -163 -88
rect -93 88 -35 100
rect -93 -88 -81 88
rect -47 -88 -35 88
rect -93 -100 -35 -88
rect 35 88 93 100
rect 35 -88 47 88
rect 81 -88 93 88
rect 35 -100 93 -88
rect 163 88 221 100
rect 163 -88 175 88
rect 209 -88 221 88
rect 163 -100 221 -88
rect 291 88 349 100
rect 291 -88 303 88
rect 337 -88 349 88
rect 291 -100 349 -88
rect 419 88 477 100
rect 419 -88 431 88
rect 465 -88 477 88
rect 419 -100 477 -88
rect 547 88 605 100
rect 547 -88 559 88
rect 593 -88 605 88
rect 547 -100 605 -88
rect 675 88 733 100
rect 675 -88 687 88
rect 721 -88 733 88
rect 675 -100 733 -88
rect 803 88 861 100
rect 803 -88 815 88
rect 849 -88 861 88
rect 803 -100 861 -88
rect 931 88 989 100
rect 931 -88 943 88
rect 977 -88 989 88
rect 931 -100 989 -88
rect 1059 88 1117 100
rect 1059 -88 1071 88
rect 1105 -88 1117 88
rect 1059 -100 1117 -88
rect 1187 88 1245 100
rect 1187 -88 1199 88
rect 1233 -88 1245 88
rect 1187 -100 1245 -88
rect 1315 88 1373 100
rect 1315 -88 1327 88
rect 1361 -88 1373 88
rect 1315 -100 1373 -88
rect 1443 88 1501 100
rect 1443 -88 1455 88
rect 1489 -88 1501 88
rect 1443 -100 1501 -88
rect 1571 88 1629 100
rect 1571 -88 1583 88
rect 1617 -88 1629 88
rect 1571 -100 1629 -88
rect 1699 88 1757 100
rect 1699 -88 1711 88
rect 1745 -88 1757 88
rect 1699 -100 1757 -88
rect 1827 88 1885 100
rect 1827 -88 1839 88
rect 1873 -88 1885 88
rect 1827 -100 1885 -88
rect 1955 88 2013 100
rect 1955 -88 1967 88
rect 2001 -88 2013 88
rect 1955 -100 2013 -88
rect 2083 88 2141 100
rect 2083 -88 2095 88
rect 2129 -88 2141 88
rect 2083 -100 2141 -88
rect 2211 88 2269 100
rect 2211 -88 2223 88
rect 2257 -88 2269 88
rect 2211 -100 2269 -88
rect 2339 88 2397 100
rect 2339 -88 2351 88
rect 2385 -88 2397 88
rect 2339 -100 2397 -88
rect 2467 88 2525 100
rect 2467 -88 2479 88
rect 2513 -88 2525 88
rect 2467 -100 2525 -88
rect 2595 88 2653 100
rect 2595 -88 2607 88
rect 2641 -88 2653 88
rect 2595 -100 2653 -88
rect 2723 88 2781 100
rect 2723 -88 2735 88
rect 2769 -88 2781 88
rect 2723 -100 2781 -88
rect 2851 88 2909 100
rect 2851 -88 2863 88
rect 2897 -88 2909 88
rect 2851 -100 2909 -88
<< pdiffc >>
rect -2897 -88 -2863 88
rect -2769 -88 -2735 88
rect -2641 -88 -2607 88
rect -2513 -88 -2479 88
rect -2385 -88 -2351 88
rect -2257 -88 -2223 88
rect -2129 -88 -2095 88
rect -2001 -88 -1967 88
rect -1873 -88 -1839 88
rect -1745 -88 -1711 88
rect -1617 -88 -1583 88
rect -1489 -88 -1455 88
rect -1361 -88 -1327 88
rect -1233 -88 -1199 88
rect -1105 -88 -1071 88
rect -977 -88 -943 88
rect -849 -88 -815 88
rect -721 -88 -687 88
rect -593 -88 -559 88
rect -465 -88 -431 88
rect -337 -88 -303 88
rect -209 -88 -175 88
rect -81 -88 -47 88
rect 47 -88 81 88
rect 175 -88 209 88
rect 303 -88 337 88
rect 431 -88 465 88
rect 559 -88 593 88
rect 687 -88 721 88
rect 815 -88 849 88
rect 943 -88 977 88
rect 1071 -88 1105 88
rect 1199 -88 1233 88
rect 1327 -88 1361 88
rect 1455 -88 1489 88
rect 1583 -88 1617 88
rect 1711 -88 1745 88
rect 1839 -88 1873 88
rect 1967 -88 2001 88
rect 2095 -88 2129 88
rect 2223 -88 2257 88
rect 2351 -88 2385 88
rect 2479 -88 2513 88
rect 2607 -88 2641 88
rect 2735 -88 2769 88
rect 2863 -88 2897 88
<< nsubdiff >>
rect -3011 249 -2915 283
rect 2915 249 3011 283
rect -3011 187 -2977 249
rect 2977 187 3011 249
rect -3011 -249 -2977 -187
rect 2977 -249 3011 -187
rect -3011 -283 -2915 -249
rect 2915 -283 3011 -249
<< nsubdiffcont >>
rect -2915 249 2915 283
rect -3011 -187 -2977 187
rect 2977 -187 3011 187
rect -2915 -283 2915 -249
<< poly >>
rect -2851 181 -2781 197
rect -2851 147 -2835 181
rect -2797 147 -2781 181
rect -2851 100 -2781 147
rect -2723 181 -2653 197
rect -2723 147 -2707 181
rect -2669 147 -2653 181
rect -2723 100 -2653 147
rect -2595 181 -2525 197
rect -2595 147 -2579 181
rect -2541 147 -2525 181
rect -2595 100 -2525 147
rect -2467 181 -2397 197
rect -2467 147 -2451 181
rect -2413 147 -2397 181
rect -2467 100 -2397 147
rect -2339 181 -2269 197
rect -2339 147 -2323 181
rect -2285 147 -2269 181
rect -2339 100 -2269 147
rect -2211 181 -2141 197
rect -2211 147 -2195 181
rect -2157 147 -2141 181
rect -2211 100 -2141 147
rect -2083 181 -2013 197
rect -2083 147 -2067 181
rect -2029 147 -2013 181
rect -2083 100 -2013 147
rect -1955 181 -1885 197
rect -1955 147 -1939 181
rect -1901 147 -1885 181
rect -1955 100 -1885 147
rect -1827 181 -1757 197
rect -1827 147 -1811 181
rect -1773 147 -1757 181
rect -1827 100 -1757 147
rect -1699 181 -1629 197
rect -1699 147 -1683 181
rect -1645 147 -1629 181
rect -1699 100 -1629 147
rect -1571 181 -1501 197
rect -1571 147 -1555 181
rect -1517 147 -1501 181
rect -1571 100 -1501 147
rect -1443 181 -1373 197
rect -1443 147 -1427 181
rect -1389 147 -1373 181
rect -1443 100 -1373 147
rect -1315 181 -1245 197
rect -1315 147 -1299 181
rect -1261 147 -1245 181
rect -1315 100 -1245 147
rect -1187 181 -1117 197
rect -1187 147 -1171 181
rect -1133 147 -1117 181
rect -1187 100 -1117 147
rect -1059 181 -989 197
rect -1059 147 -1043 181
rect -1005 147 -989 181
rect -1059 100 -989 147
rect -931 181 -861 197
rect -931 147 -915 181
rect -877 147 -861 181
rect -931 100 -861 147
rect -803 181 -733 197
rect -803 147 -787 181
rect -749 147 -733 181
rect -803 100 -733 147
rect -675 181 -605 197
rect -675 147 -659 181
rect -621 147 -605 181
rect -675 100 -605 147
rect -547 181 -477 197
rect -547 147 -531 181
rect -493 147 -477 181
rect -547 100 -477 147
rect -419 181 -349 197
rect -419 147 -403 181
rect -365 147 -349 181
rect -419 100 -349 147
rect -291 181 -221 197
rect -291 147 -275 181
rect -237 147 -221 181
rect -291 100 -221 147
rect -163 181 -93 197
rect -163 147 -147 181
rect -109 147 -93 181
rect -163 100 -93 147
rect -35 181 35 197
rect -35 147 -19 181
rect 19 147 35 181
rect -35 100 35 147
rect 93 181 163 197
rect 93 147 109 181
rect 147 147 163 181
rect 93 100 163 147
rect 221 181 291 197
rect 221 147 237 181
rect 275 147 291 181
rect 221 100 291 147
rect 349 181 419 197
rect 349 147 365 181
rect 403 147 419 181
rect 349 100 419 147
rect 477 181 547 197
rect 477 147 493 181
rect 531 147 547 181
rect 477 100 547 147
rect 605 181 675 197
rect 605 147 621 181
rect 659 147 675 181
rect 605 100 675 147
rect 733 181 803 197
rect 733 147 749 181
rect 787 147 803 181
rect 733 100 803 147
rect 861 181 931 197
rect 861 147 877 181
rect 915 147 931 181
rect 861 100 931 147
rect 989 181 1059 197
rect 989 147 1005 181
rect 1043 147 1059 181
rect 989 100 1059 147
rect 1117 181 1187 197
rect 1117 147 1133 181
rect 1171 147 1187 181
rect 1117 100 1187 147
rect 1245 181 1315 197
rect 1245 147 1261 181
rect 1299 147 1315 181
rect 1245 100 1315 147
rect 1373 181 1443 197
rect 1373 147 1389 181
rect 1427 147 1443 181
rect 1373 100 1443 147
rect 1501 181 1571 197
rect 1501 147 1517 181
rect 1555 147 1571 181
rect 1501 100 1571 147
rect 1629 181 1699 197
rect 1629 147 1645 181
rect 1683 147 1699 181
rect 1629 100 1699 147
rect 1757 181 1827 197
rect 1757 147 1773 181
rect 1811 147 1827 181
rect 1757 100 1827 147
rect 1885 181 1955 197
rect 1885 147 1901 181
rect 1939 147 1955 181
rect 1885 100 1955 147
rect 2013 181 2083 197
rect 2013 147 2029 181
rect 2067 147 2083 181
rect 2013 100 2083 147
rect 2141 181 2211 197
rect 2141 147 2157 181
rect 2195 147 2211 181
rect 2141 100 2211 147
rect 2269 181 2339 197
rect 2269 147 2285 181
rect 2323 147 2339 181
rect 2269 100 2339 147
rect 2397 181 2467 197
rect 2397 147 2413 181
rect 2451 147 2467 181
rect 2397 100 2467 147
rect 2525 181 2595 197
rect 2525 147 2541 181
rect 2579 147 2595 181
rect 2525 100 2595 147
rect 2653 181 2723 197
rect 2653 147 2669 181
rect 2707 147 2723 181
rect 2653 100 2723 147
rect 2781 181 2851 197
rect 2781 147 2797 181
rect 2835 147 2851 181
rect 2781 100 2851 147
rect -2851 -147 -2781 -100
rect -2851 -181 -2835 -147
rect -2797 -181 -2781 -147
rect -2851 -197 -2781 -181
rect -2723 -147 -2653 -100
rect -2723 -181 -2707 -147
rect -2669 -181 -2653 -147
rect -2723 -197 -2653 -181
rect -2595 -147 -2525 -100
rect -2595 -181 -2579 -147
rect -2541 -181 -2525 -147
rect -2595 -197 -2525 -181
rect -2467 -147 -2397 -100
rect -2467 -181 -2451 -147
rect -2413 -181 -2397 -147
rect -2467 -197 -2397 -181
rect -2339 -147 -2269 -100
rect -2339 -181 -2323 -147
rect -2285 -181 -2269 -147
rect -2339 -197 -2269 -181
rect -2211 -147 -2141 -100
rect -2211 -181 -2195 -147
rect -2157 -181 -2141 -147
rect -2211 -197 -2141 -181
rect -2083 -147 -2013 -100
rect -2083 -181 -2067 -147
rect -2029 -181 -2013 -147
rect -2083 -197 -2013 -181
rect -1955 -147 -1885 -100
rect -1955 -181 -1939 -147
rect -1901 -181 -1885 -147
rect -1955 -197 -1885 -181
rect -1827 -147 -1757 -100
rect -1827 -181 -1811 -147
rect -1773 -181 -1757 -147
rect -1827 -197 -1757 -181
rect -1699 -147 -1629 -100
rect -1699 -181 -1683 -147
rect -1645 -181 -1629 -147
rect -1699 -197 -1629 -181
rect -1571 -147 -1501 -100
rect -1571 -181 -1555 -147
rect -1517 -181 -1501 -147
rect -1571 -197 -1501 -181
rect -1443 -147 -1373 -100
rect -1443 -181 -1427 -147
rect -1389 -181 -1373 -147
rect -1443 -197 -1373 -181
rect -1315 -147 -1245 -100
rect -1315 -181 -1299 -147
rect -1261 -181 -1245 -147
rect -1315 -197 -1245 -181
rect -1187 -147 -1117 -100
rect -1187 -181 -1171 -147
rect -1133 -181 -1117 -147
rect -1187 -197 -1117 -181
rect -1059 -147 -989 -100
rect -1059 -181 -1043 -147
rect -1005 -181 -989 -147
rect -1059 -197 -989 -181
rect -931 -147 -861 -100
rect -931 -181 -915 -147
rect -877 -181 -861 -147
rect -931 -197 -861 -181
rect -803 -147 -733 -100
rect -803 -181 -787 -147
rect -749 -181 -733 -147
rect -803 -197 -733 -181
rect -675 -147 -605 -100
rect -675 -181 -659 -147
rect -621 -181 -605 -147
rect -675 -197 -605 -181
rect -547 -147 -477 -100
rect -547 -181 -531 -147
rect -493 -181 -477 -147
rect -547 -197 -477 -181
rect -419 -147 -349 -100
rect -419 -181 -403 -147
rect -365 -181 -349 -147
rect -419 -197 -349 -181
rect -291 -147 -221 -100
rect -291 -181 -275 -147
rect -237 -181 -221 -147
rect -291 -197 -221 -181
rect -163 -147 -93 -100
rect -163 -181 -147 -147
rect -109 -181 -93 -147
rect -163 -197 -93 -181
rect -35 -147 35 -100
rect -35 -181 -19 -147
rect 19 -181 35 -147
rect -35 -197 35 -181
rect 93 -147 163 -100
rect 93 -181 109 -147
rect 147 -181 163 -147
rect 93 -197 163 -181
rect 221 -147 291 -100
rect 221 -181 237 -147
rect 275 -181 291 -147
rect 221 -197 291 -181
rect 349 -147 419 -100
rect 349 -181 365 -147
rect 403 -181 419 -147
rect 349 -197 419 -181
rect 477 -147 547 -100
rect 477 -181 493 -147
rect 531 -181 547 -147
rect 477 -197 547 -181
rect 605 -147 675 -100
rect 605 -181 621 -147
rect 659 -181 675 -147
rect 605 -197 675 -181
rect 733 -147 803 -100
rect 733 -181 749 -147
rect 787 -181 803 -147
rect 733 -197 803 -181
rect 861 -147 931 -100
rect 861 -181 877 -147
rect 915 -181 931 -147
rect 861 -197 931 -181
rect 989 -147 1059 -100
rect 989 -181 1005 -147
rect 1043 -181 1059 -147
rect 989 -197 1059 -181
rect 1117 -147 1187 -100
rect 1117 -181 1133 -147
rect 1171 -181 1187 -147
rect 1117 -197 1187 -181
rect 1245 -147 1315 -100
rect 1245 -181 1261 -147
rect 1299 -181 1315 -147
rect 1245 -197 1315 -181
rect 1373 -147 1443 -100
rect 1373 -181 1389 -147
rect 1427 -181 1443 -147
rect 1373 -197 1443 -181
rect 1501 -147 1571 -100
rect 1501 -181 1517 -147
rect 1555 -181 1571 -147
rect 1501 -197 1571 -181
rect 1629 -147 1699 -100
rect 1629 -181 1645 -147
rect 1683 -181 1699 -147
rect 1629 -197 1699 -181
rect 1757 -147 1827 -100
rect 1757 -181 1773 -147
rect 1811 -181 1827 -147
rect 1757 -197 1827 -181
rect 1885 -147 1955 -100
rect 1885 -181 1901 -147
rect 1939 -181 1955 -147
rect 1885 -197 1955 -181
rect 2013 -147 2083 -100
rect 2013 -181 2029 -147
rect 2067 -181 2083 -147
rect 2013 -197 2083 -181
rect 2141 -147 2211 -100
rect 2141 -181 2157 -147
rect 2195 -181 2211 -147
rect 2141 -197 2211 -181
rect 2269 -147 2339 -100
rect 2269 -181 2285 -147
rect 2323 -181 2339 -147
rect 2269 -197 2339 -181
rect 2397 -147 2467 -100
rect 2397 -181 2413 -147
rect 2451 -181 2467 -147
rect 2397 -197 2467 -181
rect 2525 -147 2595 -100
rect 2525 -181 2541 -147
rect 2579 -181 2595 -147
rect 2525 -197 2595 -181
rect 2653 -147 2723 -100
rect 2653 -181 2669 -147
rect 2707 -181 2723 -147
rect 2653 -197 2723 -181
rect 2781 -147 2851 -100
rect 2781 -181 2797 -147
rect 2835 -181 2851 -147
rect 2781 -197 2851 -181
<< polycont >>
rect -2835 147 -2797 181
rect -2707 147 -2669 181
rect -2579 147 -2541 181
rect -2451 147 -2413 181
rect -2323 147 -2285 181
rect -2195 147 -2157 181
rect -2067 147 -2029 181
rect -1939 147 -1901 181
rect -1811 147 -1773 181
rect -1683 147 -1645 181
rect -1555 147 -1517 181
rect -1427 147 -1389 181
rect -1299 147 -1261 181
rect -1171 147 -1133 181
rect -1043 147 -1005 181
rect -915 147 -877 181
rect -787 147 -749 181
rect -659 147 -621 181
rect -531 147 -493 181
rect -403 147 -365 181
rect -275 147 -237 181
rect -147 147 -109 181
rect -19 147 19 181
rect 109 147 147 181
rect 237 147 275 181
rect 365 147 403 181
rect 493 147 531 181
rect 621 147 659 181
rect 749 147 787 181
rect 877 147 915 181
rect 1005 147 1043 181
rect 1133 147 1171 181
rect 1261 147 1299 181
rect 1389 147 1427 181
rect 1517 147 1555 181
rect 1645 147 1683 181
rect 1773 147 1811 181
rect 1901 147 1939 181
rect 2029 147 2067 181
rect 2157 147 2195 181
rect 2285 147 2323 181
rect 2413 147 2451 181
rect 2541 147 2579 181
rect 2669 147 2707 181
rect 2797 147 2835 181
rect -2835 -181 -2797 -147
rect -2707 -181 -2669 -147
rect -2579 -181 -2541 -147
rect -2451 -181 -2413 -147
rect -2323 -181 -2285 -147
rect -2195 -181 -2157 -147
rect -2067 -181 -2029 -147
rect -1939 -181 -1901 -147
rect -1811 -181 -1773 -147
rect -1683 -181 -1645 -147
rect -1555 -181 -1517 -147
rect -1427 -181 -1389 -147
rect -1299 -181 -1261 -147
rect -1171 -181 -1133 -147
rect -1043 -181 -1005 -147
rect -915 -181 -877 -147
rect -787 -181 -749 -147
rect -659 -181 -621 -147
rect -531 -181 -493 -147
rect -403 -181 -365 -147
rect -275 -181 -237 -147
rect -147 -181 -109 -147
rect -19 -181 19 -147
rect 109 -181 147 -147
rect 237 -181 275 -147
rect 365 -181 403 -147
rect 493 -181 531 -147
rect 621 -181 659 -147
rect 749 -181 787 -147
rect 877 -181 915 -147
rect 1005 -181 1043 -147
rect 1133 -181 1171 -147
rect 1261 -181 1299 -147
rect 1389 -181 1427 -147
rect 1517 -181 1555 -147
rect 1645 -181 1683 -147
rect 1773 -181 1811 -147
rect 1901 -181 1939 -147
rect 2029 -181 2067 -147
rect 2157 -181 2195 -147
rect 2285 -181 2323 -147
rect 2413 -181 2451 -147
rect 2541 -181 2579 -147
rect 2669 -181 2707 -147
rect 2797 -181 2835 -147
<< locali >>
rect -3011 249 -2915 283
rect 2915 249 3011 283
rect -3011 187 -2977 249
rect 2977 187 3011 249
rect -2851 147 -2835 181
rect -2797 147 -2781 181
rect -2723 147 -2707 181
rect -2669 147 -2653 181
rect -2595 147 -2579 181
rect -2541 147 -2525 181
rect -2467 147 -2451 181
rect -2413 147 -2397 181
rect -2339 147 -2323 181
rect -2285 147 -2269 181
rect -2211 147 -2195 181
rect -2157 147 -2141 181
rect -2083 147 -2067 181
rect -2029 147 -2013 181
rect -1955 147 -1939 181
rect -1901 147 -1885 181
rect -1827 147 -1811 181
rect -1773 147 -1757 181
rect -1699 147 -1683 181
rect -1645 147 -1629 181
rect -1571 147 -1555 181
rect -1517 147 -1501 181
rect -1443 147 -1427 181
rect -1389 147 -1373 181
rect -1315 147 -1299 181
rect -1261 147 -1245 181
rect -1187 147 -1171 181
rect -1133 147 -1117 181
rect -1059 147 -1043 181
rect -1005 147 -989 181
rect -931 147 -915 181
rect -877 147 -861 181
rect -803 147 -787 181
rect -749 147 -733 181
rect -675 147 -659 181
rect -621 147 -605 181
rect -547 147 -531 181
rect -493 147 -477 181
rect -419 147 -403 181
rect -365 147 -349 181
rect -291 147 -275 181
rect -237 147 -221 181
rect -163 147 -147 181
rect -109 147 -93 181
rect -35 147 -19 181
rect 19 147 35 181
rect 93 147 109 181
rect 147 147 163 181
rect 221 147 237 181
rect 275 147 291 181
rect 349 147 365 181
rect 403 147 419 181
rect 477 147 493 181
rect 531 147 547 181
rect 605 147 621 181
rect 659 147 675 181
rect 733 147 749 181
rect 787 147 803 181
rect 861 147 877 181
rect 915 147 931 181
rect 989 147 1005 181
rect 1043 147 1059 181
rect 1117 147 1133 181
rect 1171 147 1187 181
rect 1245 147 1261 181
rect 1299 147 1315 181
rect 1373 147 1389 181
rect 1427 147 1443 181
rect 1501 147 1517 181
rect 1555 147 1571 181
rect 1629 147 1645 181
rect 1683 147 1699 181
rect 1757 147 1773 181
rect 1811 147 1827 181
rect 1885 147 1901 181
rect 1939 147 1955 181
rect 2013 147 2029 181
rect 2067 147 2083 181
rect 2141 147 2157 181
rect 2195 147 2211 181
rect 2269 147 2285 181
rect 2323 147 2339 181
rect 2397 147 2413 181
rect 2451 147 2467 181
rect 2525 147 2541 181
rect 2579 147 2595 181
rect 2653 147 2669 181
rect 2707 147 2723 181
rect 2781 147 2797 181
rect 2835 147 2851 181
rect -2897 88 -2863 104
rect -2897 -104 -2863 -88
rect -2769 88 -2735 104
rect -2769 -104 -2735 -88
rect -2641 88 -2607 104
rect -2641 -104 -2607 -88
rect -2513 88 -2479 104
rect -2513 -104 -2479 -88
rect -2385 88 -2351 104
rect -2385 -104 -2351 -88
rect -2257 88 -2223 104
rect -2257 -104 -2223 -88
rect -2129 88 -2095 104
rect -2129 -104 -2095 -88
rect -2001 88 -1967 104
rect -2001 -104 -1967 -88
rect -1873 88 -1839 104
rect -1873 -104 -1839 -88
rect -1745 88 -1711 104
rect -1745 -104 -1711 -88
rect -1617 88 -1583 104
rect -1617 -104 -1583 -88
rect -1489 88 -1455 104
rect -1489 -104 -1455 -88
rect -1361 88 -1327 104
rect -1361 -104 -1327 -88
rect -1233 88 -1199 104
rect -1233 -104 -1199 -88
rect -1105 88 -1071 104
rect -1105 -104 -1071 -88
rect -977 88 -943 104
rect -977 -104 -943 -88
rect -849 88 -815 104
rect -849 -104 -815 -88
rect -721 88 -687 104
rect -721 -104 -687 -88
rect -593 88 -559 104
rect -593 -104 -559 -88
rect -465 88 -431 104
rect -465 -104 -431 -88
rect -337 88 -303 104
rect -337 -104 -303 -88
rect -209 88 -175 104
rect -209 -104 -175 -88
rect -81 88 -47 104
rect -81 -104 -47 -88
rect 47 88 81 104
rect 47 -104 81 -88
rect 175 88 209 104
rect 175 -104 209 -88
rect 303 88 337 104
rect 303 -104 337 -88
rect 431 88 465 104
rect 431 -104 465 -88
rect 559 88 593 104
rect 559 -104 593 -88
rect 687 88 721 104
rect 687 -104 721 -88
rect 815 88 849 104
rect 815 -104 849 -88
rect 943 88 977 104
rect 943 -104 977 -88
rect 1071 88 1105 104
rect 1071 -104 1105 -88
rect 1199 88 1233 104
rect 1199 -104 1233 -88
rect 1327 88 1361 104
rect 1327 -104 1361 -88
rect 1455 88 1489 104
rect 1455 -104 1489 -88
rect 1583 88 1617 104
rect 1583 -104 1617 -88
rect 1711 88 1745 104
rect 1711 -104 1745 -88
rect 1839 88 1873 104
rect 1839 -104 1873 -88
rect 1967 88 2001 104
rect 1967 -104 2001 -88
rect 2095 88 2129 104
rect 2095 -104 2129 -88
rect 2223 88 2257 104
rect 2223 -104 2257 -88
rect 2351 88 2385 104
rect 2351 -104 2385 -88
rect 2479 88 2513 104
rect 2479 -104 2513 -88
rect 2607 88 2641 104
rect 2607 -104 2641 -88
rect 2735 88 2769 104
rect 2735 -104 2769 -88
rect 2863 88 2897 104
rect 2863 -104 2897 -88
rect -2851 -181 -2835 -147
rect -2797 -181 -2781 -147
rect -2723 -181 -2707 -147
rect -2669 -181 -2653 -147
rect -2595 -181 -2579 -147
rect -2541 -181 -2525 -147
rect -2467 -181 -2451 -147
rect -2413 -181 -2397 -147
rect -2339 -181 -2323 -147
rect -2285 -181 -2269 -147
rect -2211 -181 -2195 -147
rect -2157 -181 -2141 -147
rect -2083 -181 -2067 -147
rect -2029 -181 -2013 -147
rect -1955 -181 -1939 -147
rect -1901 -181 -1885 -147
rect -1827 -181 -1811 -147
rect -1773 -181 -1757 -147
rect -1699 -181 -1683 -147
rect -1645 -181 -1629 -147
rect -1571 -181 -1555 -147
rect -1517 -181 -1501 -147
rect -1443 -181 -1427 -147
rect -1389 -181 -1373 -147
rect -1315 -181 -1299 -147
rect -1261 -181 -1245 -147
rect -1187 -181 -1171 -147
rect -1133 -181 -1117 -147
rect -1059 -181 -1043 -147
rect -1005 -181 -989 -147
rect -931 -181 -915 -147
rect -877 -181 -861 -147
rect -803 -181 -787 -147
rect -749 -181 -733 -147
rect -675 -181 -659 -147
rect -621 -181 -605 -147
rect -547 -181 -531 -147
rect -493 -181 -477 -147
rect -419 -181 -403 -147
rect -365 -181 -349 -147
rect -291 -181 -275 -147
rect -237 -181 -221 -147
rect -163 -181 -147 -147
rect -109 -181 -93 -147
rect -35 -181 -19 -147
rect 19 -181 35 -147
rect 93 -181 109 -147
rect 147 -181 163 -147
rect 221 -181 237 -147
rect 275 -181 291 -147
rect 349 -181 365 -147
rect 403 -181 419 -147
rect 477 -181 493 -147
rect 531 -181 547 -147
rect 605 -181 621 -147
rect 659 -181 675 -147
rect 733 -181 749 -147
rect 787 -181 803 -147
rect 861 -181 877 -147
rect 915 -181 931 -147
rect 989 -181 1005 -147
rect 1043 -181 1059 -147
rect 1117 -181 1133 -147
rect 1171 -181 1187 -147
rect 1245 -181 1261 -147
rect 1299 -181 1315 -147
rect 1373 -181 1389 -147
rect 1427 -181 1443 -147
rect 1501 -181 1517 -147
rect 1555 -181 1571 -147
rect 1629 -181 1645 -147
rect 1683 -181 1699 -147
rect 1757 -181 1773 -147
rect 1811 -181 1827 -147
rect 1885 -181 1901 -147
rect 1939 -181 1955 -147
rect 2013 -181 2029 -147
rect 2067 -181 2083 -147
rect 2141 -181 2157 -147
rect 2195 -181 2211 -147
rect 2269 -181 2285 -147
rect 2323 -181 2339 -147
rect 2397 -181 2413 -147
rect 2451 -181 2467 -147
rect 2525 -181 2541 -147
rect 2579 -181 2595 -147
rect 2653 -181 2669 -147
rect 2707 -181 2723 -147
rect 2781 -181 2797 -147
rect 2835 -181 2851 -147
rect -3011 -249 -2977 -187
rect 2977 -249 3011 -187
rect -3011 -283 -2915 -249
rect 2915 -283 3011 -249
<< viali >>
rect -2835 147 -2797 181
rect -2707 147 -2669 181
rect -2579 147 -2541 181
rect -2451 147 -2413 181
rect -2323 147 -2285 181
rect -2195 147 -2157 181
rect -2067 147 -2029 181
rect -1939 147 -1901 181
rect -1811 147 -1773 181
rect -1683 147 -1645 181
rect -1555 147 -1517 181
rect -1427 147 -1389 181
rect -1299 147 -1261 181
rect -1171 147 -1133 181
rect -1043 147 -1005 181
rect -915 147 -877 181
rect -787 147 -749 181
rect -659 147 -621 181
rect -531 147 -493 181
rect -403 147 -365 181
rect -275 147 -237 181
rect -147 147 -109 181
rect -19 147 19 181
rect 109 147 147 181
rect 237 147 275 181
rect 365 147 403 181
rect 493 147 531 181
rect 621 147 659 181
rect 749 147 787 181
rect 877 147 915 181
rect 1005 147 1043 181
rect 1133 147 1171 181
rect 1261 147 1299 181
rect 1389 147 1427 181
rect 1517 147 1555 181
rect 1645 147 1683 181
rect 1773 147 1811 181
rect 1901 147 1939 181
rect 2029 147 2067 181
rect 2157 147 2195 181
rect 2285 147 2323 181
rect 2413 147 2451 181
rect 2541 147 2579 181
rect 2669 147 2707 181
rect 2797 147 2835 181
rect -2897 -88 -2863 88
rect -2769 -88 -2735 88
rect -2641 -88 -2607 88
rect -2513 -88 -2479 88
rect -2385 -88 -2351 88
rect -2257 -88 -2223 88
rect -2129 -88 -2095 88
rect -2001 -88 -1967 88
rect -1873 -88 -1839 88
rect -1745 -88 -1711 88
rect -1617 -88 -1583 88
rect -1489 -88 -1455 88
rect -1361 -88 -1327 88
rect -1233 -88 -1199 88
rect -1105 -88 -1071 88
rect -977 -88 -943 88
rect -849 -88 -815 88
rect -721 -88 -687 88
rect -593 -88 -559 88
rect -465 -88 -431 88
rect -337 -88 -303 88
rect -209 -88 -175 88
rect -81 -88 -47 88
rect 47 -88 81 88
rect 175 -88 209 88
rect 303 -88 337 88
rect 431 -88 465 88
rect 559 -88 593 88
rect 687 -88 721 88
rect 815 -88 849 88
rect 943 -88 977 88
rect 1071 -88 1105 88
rect 1199 -88 1233 88
rect 1327 -88 1361 88
rect 1455 -88 1489 88
rect 1583 -88 1617 88
rect 1711 -88 1745 88
rect 1839 -88 1873 88
rect 1967 -88 2001 88
rect 2095 -88 2129 88
rect 2223 -88 2257 88
rect 2351 -88 2385 88
rect 2479 -88 2513 88
rect 2607 -88 2641 88
rect 2735 -88 2769 88
rect 2863 -88 2897 88
rect -2835 -181 -2797 -147
rect -2707 -181 -2669 -147
rect -2579 -181 -2541 -147
rect -2451 -181 -2413 -147
rect -2323 -181 -2285 -147
rect -2195 -181 -2157 -147
rect -2067 -181 -2029 -147
rect -1939 -181 -1901 -147
rect -1811 -181 -1773 -147
rect -1683 -181 -1645 -147
rect -1555 -181 -1517 -147
rect -1427 -181 -1389 -147
rect -1299 -181 -1261 -147
rect -1171 -181 -1133 -147
rect -1043 -181 -1005 -147
rect -915 -181 -877 -147
rect -787 -181 -749 -147
rect -659 -181 -621 -147
rect -531 -181 -493 -147
rect -403 -181 -365 -147
rect -275 -181 -237 -147
rect -147 -181 -109 -147
rect -19 -181 19 -147
rect 109 -181 147 -147
rect 237 -181 275 -147
rect 365 -181 403 -147
rect 493 -181 531 -147
rect 621 -181 659 -147
rect 749 -181 787 -147
rect 877 -181 915 -147
rect 1005 -181 1043 -147
rect 1133 -181 1171 -147
rect 1261 -181 1299 -147
rect 1389 -181 1427 -147
rect 1517 -181 1555 -147
rect 1645 -181 1683 -147
rect 1773 -181 1811 -147
rect 1901 -181 1939 -147
rect 2029 -181 2067 -147
rect 2157 -181 2195 -147
rect 2285 -181 2323 -147
rect 2413 -181 2451 -147
rect 2541 -181 2579 -147
rect 2669 -181 2707 -147
rect 2797 -181 2835 -147
<< metal1 >>
rect -2847 181 -2785 187
rect -2847 147 -2835 181
rect -2797 147 -2785 181
rect -2847 141 -2785 147
rect -2719 181 -2657 187
rect -2719 147 -2707 181
rect -2669 147 -2657 181
rect -2719 141 -2657 147
rect -2591 181 -2529 187
rect -2591 147 -2579 181
rect -2541 147 -2529 181
rect -2591 141 -2529 147
rect -2463 181 -2401 187
rect -2463 147 -2451 181
rect -2413 147 -2401 181
rect -2463 141 -2401 147
rect -2335 181 -2273 187
rect -2335 147 -2323 181
rect -2285 147 -2273 181
rect -2335 141 -2273 147
rect -2207 181 -2145 187
rect -2207 147 -2195 181
rect -2157 147 -2145 181
rect -2207 141 -2145 147
rect -2079 181 -2017 187
rect -2079 147 -2067 181
rect -2029 147 -2017 181
rect -2079 141 -2017 147
rect -1951 181 -1889 187
rect -1951 147 -1939 181
rect -1901 147 -1889 181
rect -1951 141 -1889 147
rect -1823 181 -1761 187
rect -1823 147 -1811 181
rect -1773 147 -1761 181
rect -1823 141 -1761 147
rect -1695 181 -1633 187
rect -1695 147 -1683 181
rect -1645 147 -1633 181
rect -1695 141 -1633 147
rect -1567 181 -1505 187
rect -1567 147 -1555 181
rect -1517 147 -1505 181
rect -1567 141 -1505 147
rect -1439 181 -1377 187
rect -1439 147 -1427 181
rect -1389 147 -1377 181
rect -1439 141 -1377 147
rect -1311 181 -1249 187
rect -1311 147 -1299 181
rect -1261 147 -1249 181
rect -1311 141 -1249 147
rect -1183 181 -1121 187
rect -1183 147 -1171 181
rect -1133 147 -1121 181
rect -1183 141 -1121 147
rect -1055 181 -993 187
rect -1055 147 -1043 181
rect -1005 147 -993 181
rect -1055 141 -993 147
rect -927 181 -865 187
rect -927 147 -915 181
rect -877 147 -865 181
rect -927 141 -865 147
rect -799 181 -737 187
rect -799 147 -787 181
rect -749 147 -737 181
rect -799 141 -737 147
rect -671 181 -609 187
rect -671 147 -659 181
rect -621 147 -609 181
rect -671 141 -609 147
rect -543 181 -481 187
rect -543 147 -531 181
rect -493 147 -481 181
rect -543 141 -481 147
rect -415 181 -353 187
rect -415 147 -403 181
rect -365 147 -353 181
rect -415 141 -353 147
rect -287 181 -225 187
rect -287 147 -275 181
rect -237 147 -225 181
rect -287 141 -225 147
rect -159 181 -97 187
rect -159 147 -147 181
rect -109 147 -97 181
rect -159 141 -97 147
rect -31 181 31 187
rect -31 147 -19 181
rect 19 147 31 181
rect -31 141 31 147
rect 97 181 159 187
rect 97 147 109 181
rect 147 147 159 181
rect 97 141 159 147
rect 225 181 287 187
rect 225 147 237 181
rect 275 147 287 181
rect 225 141 287 147
rect 353 181 415 187
rect 353 147 365 181
rect 403 147 415 181
rect 353 141 415 147
rect 481 181 543 187
rect 481 147 493 181
rect 531 147 543 181
rect 481 141 543 147
rect 609 181 671 187
rect 609 147 621 181
rect 659 147 671 181
rect 609 141 671 147
rect 737 181 799 187
rect 737 147 749 181
rect 787 147 799 181
rect 737 141 799 147
rect 865 181 927 187
rect 865 147 877 181
rect 915 147 927 181
rect 865 141 927 147
rect 993 181 1055 187
rect 993 147 1005 181
rect 1043 147 1055 181
rect 993 141 1055 147
rect 1121 181 1183 187
rect 1121 147 1133 181
rect 1171 147 1183 181
rect 1121 141 1183 147
rect 1249 181 1311 187
rect 1249 147 1261 181
rect 1299 147 1311 181
rect 1249 141 1311 147
rect 1377 181 1439 187
rect 1377 147 1389 181
rect 1427 147 1439 181
rect 1377 141 1439 147
rect 1505 181 1567 187
rect 1505 147 1517 181
rect 1555 147 1567 181
rect 1505 141 1567 147
rect 1633 181 1695 187
rect 1633 147 1645 181
rect 1683 147 1695 181
rect 1633 141 1695 147
rect 1761 181 1823 187
rect 1761 147 1773 181
rect 1811 147 1823 181
rect 1761 141 1823 147
rect 1889 181 1951 187
rect 1889 147 1901 181
rect 1939 147 1951 181
rect 1889 141 1951 147
rect 2017 181 2079 187
rect 2017 147 2029 181
rect 2067 147 2079 181
rect 2017 141 2079 147
rect 2145 181 2207 187
rect 2145 147 2157 181
rect 2195 147 2207 181
rect 2145 141 2207 147
rect 2273 181 2335 187
rect 2273 147 2285 181
rect 2323 147 2335 181
rect 2273 141 2335 147
rect 2401 181 2463 187
rect 2401 147 2413 181
rect 2451 147 2463 181
rect 2401 141 2463 147
rect 2529 181 2591 187
rect 2529 147 2541 181
rect 2579 147 2591 181
rect 2529 141 2591 147
rect 2657 181 2719 187
rect 2657 147 2669 181
rect 2707 147 2719 181
rect 2657 141 2719 147
rect 2785 181 2847 187
rect 2785 147 2797 181
rect 2835 147 2847 181
rect 2785 141 2847 147
rect -2903 88 -2857 100
rect -2903 -88 -2897 88
rect -2863 -88 -2857 88
rect -2903 -100 -2857 -88
rect -2775 88 -2729 100
rect -2775 -88 -2769 88
rect -2735 -88 -2729 88
rect -2775 -100 -2729 -88
rect -2647 88 -2601 100
rect -2647 -88 -2641 88
rect -2607 -88 -2601 88
rect -2647 -100 -2601 -88
rect -2519 88 -2473 100
rect -2519 -88 -2513 88
rect -2479 -88 -2473 88
rect -2519 -100 -2473 -88
rect -2391 88 -2345 100
rect -2391 -88 -2385 88
rect -2351 -88 -2345 88
rect -2391 -100 -2345 -88
rect -2263 88 -2217 100
rect -2263 -88 -2257 88
rect -2223 -88 -2217 88
rect -2263 -100 -2217 -88
rect -2135 88 -2089 100
rect -2135 -88 -2129 88
rect -2095 -88 -2089 88
rect -2135 -100 -2089 -88
rect -2007 88 -1961 100
rect -2007 -88 -2001 88
rect -1967 -88 -1961 88
rect -2007 -100 -1961 -88
rect -1879 88 -1833 100
rect -1879 -88 -1873 88
rect -1839 -88 -1833 88
rect -1879 -100 -1833 -88
rect -1751 88 -1705 100
rect -1751 -88 -1745 88
rect -1711 -88 -1705 88
rect -1751 -100 -1705 -88
rect -1623 88 -1577 100
rect -1623 -88 -1617 88
rect -1583 -88 -1577 88
rect -1623 -100 -1577 -88
rect -1495 88 -1449 100
rect -1495 -88 -1489 88
rect -1455 -88 -1449 88
rect -1495 -100 -1449 -88
rect -1367 88 -1321 100
rect -1367 -88 -1361 88
rect -1327 -88 -1321 88
rect -1367 -100 -1321 -88
rect -1239 88 -1193 100
rect -1239 -88 -1233 88
rect -1199 -88 -1193 88
rect -1239 -100 -1193 -88
rect -1111 88 -1065 100
rect -1111 -88 -1105 88
rect -1071 -88 -1065 88
rect -1111 -100 -1065 -88
rect -983 88 -937 100
rect -983 -88 -977 88
rect -943 -88 -937 88
rect -983 -100 -937 -88
rect -855 88 -809 100
rect -855 -88 -849 88
rect -815 -88 -809 88
rect -855 -100 -809 -88
rect -727 88 -681 100
rect -727 -88 -721 88
rect -687 -88 -681 88
rect -727 -100 -681 -88
rect -599 88 -553 100
rect -599 -88 -593 88
rect -559 -88 -553 88
rect -599 -100 -553 -88
rect -471 88 -425 100
rect -471 -88 -465 88
rect -431 -88 -425 88
rect -471 -100 -425 -88
rect -343 88 -297 100
rect -343 -88 -337 88
rect -303 -88 -297 88
rect -343 -100 -297 -88
rect -215 88 -169 100
rect -215 -88 -209 88
rect -175 -88 -169 88
rect -215 -100 -169 -88
rect -87 88 -41 100
rect -87 -88 -81 88
rect -47 -88 -41 88
rect -87 -100 -41 -88
rect 41 88 87 100
rect 41 -88 47 88
rect 81 -88 87 88
rect 41 -100 87 -88
rect 169 88 215 100
rect 169 -88 175 88
rect 209 -88 215 88
rect 169 -100 215 -88
rect 297 88 343 100
rect 297 -88 303 88
rect 337 -88 343 88
rect 297 -100 343 -88
rect 425 88 471 100
rect 425 -88 431 88
rect 465 -88 471 88
rect 425 -100 471 -88
rect 553 88 599 100
rect 553 -88 559 88
rect 593 -88 599 88
rect 553 -100 599 -88
rect 681 88 727 100
rect 681 -88 687 88
rect 721 -88 727 88
rect 681 -100 727 -88
rect 809 88 855 100
rect 809 -88 815 88
rect 849 -88 855 88
rect 809 -100 855 -88
rect 937 88 983 100
rect 937 -88 943 88
rect 977 -88 983 88
rect 937 -100 983 -88
rect 1065 88 1111 100
rect 1065 -88 1071 88
rect 1105 -88 1111 88
rect 1065 -100 1111 -88
rect 1193 88 1239 100
rect 1193 -88 1199 88
rect 1233 -88 1239 88
rect 1193 -100 1239 -88
rect 1321 88 1367 100
rect 1321 -88 1327 88
rect 1361 -88 1367 88
rect 1321 -100 1367 -88
rect 1449 88 1495 100
rect 1449 -88 1455 88
rect 1489 -88 1495 88
rect 1449 -100 1495 -88
rect 1577 88 1623 100
rect 1577 -88 1583 88
rect 1617 -88 1623 88
rect 1577 -100 1623 -88
rect 1705 88 1751 100
rect 1705 -88 1711 88
rect 1745 -88 1751 88
rect 1705 -100 1751 -88
rect 1833 88 1879 100
rect 1833 -88 1839 88
rect 1873 -88 1879 88
rect 1833 -100 1879 -88
rect 1961 88 2007 100
rect 1961 -88 1967 88
rect 2001 -88 2007 88
rect 1961 -100 2007 -88
rect 2089 88 2135 100
rect 2089 -88 2095 88
rect 2129 -88 2135 88
rect 2089 -100 2135 -88
rect 2217 88 2263 100
rect 2217 -88 2223 88
rect 2257 -88 2263 88
rect 2217 -100 2263 -88
rect 2345 88 2391 100
rect 2345 -88 2351 88
rect 2385 -88 2391 88
rect 2345 -100 2391 -88
rect 2473 88 2519 100
rect 2473 -88 2479 88
rect 2513 -88 2519 88
rect 2473 -100 2519 -88
rect 2601 88 2647 100
rect 2601 -88 2607 88
rect 2641 -88 2647 88
rect 2601 -100 2647 -88
rect 2729 88 2775 100
rect 2729 -88 2735 88
rect 2769 -88 2775 88
rect 2729 -100 2775 -88
rect 2857 88 2903 100
rect 2857 -88 2863 88
rect 2897 -88 2903 88
rect 2857 -100 2903 -88
rect -2847 -147 -2785 -141
rect -2847 -181 -2835 -147
rect -2797 -181 -2785 -147
rect -2847 -187 -2785 -181
rect -2719 -147 -2657 -141
rect -2719 -181 -2707 -147
rect -2669 -181 -2657 -147
rect -2719 -187 -2657 -181
rect -2591 -147 -2529 -141
rect -2591 -181 -2579 -147
rect -2541 -181 -2529 -147
rect -2591 -187 -2529 -181
rect -2463 -147 -2401 -141
rect -2463 -181 -2451 -147
rect -2413 -181 -2401 -147
rect -2463 -187 -2401 -181
rect -2335 -147 -2273 -141
rect -2335 -181 -2323 -147
rect -2285 -181 -2273 -147
rect -2335 -187 -2273 -181
rect -2207 -147 -2145 -141
rect -2207 -181 -2195 -147
rect -2157 -181 -2145 -147
rect -2207 -187 -2145 -181
rect -2079 -147 -2017 -141
rect -2079 -181 -2067 -147
rect -2029 -181 -2017 -147
rect -2079 -187 -2017 -181
rect -1951 -147 -1889 -141
rect -1951 -181 -1939 -147
rect -1901 -181 -1889 -147
rect -1951 -187 -1889 -181
rect -1823 -147 -1761 -141
rect -1823 -181 -1811 -147
rect -1773 -181 -1761 -147
rect -1823 -187 -1761 -181
rect -1695 -147 -1633 -141
rect -1695 -181 -1683 -147
rect -1645 -181 -1633 -147
rect -1695 -187 -1633 -181
rect -1567 -147 -1505 -141
rect -1567 -181 -1555 -147
rect -1517 -181 -1505 -147
rect -1567 -187 -1505 -181
rect -1439 -147 -1377 -141
rect -1439 -181 -1427 -147
rect -1389 -181 -1377 -147
rect -1439 -187 -1377 -181
rect -1311 -147 -1249 -141
rect -1311 -181 -1299 -147
rect -1261 -181 -1249 -147
rect -1311 -187 -1249 -181
rect -1183 -147 -1121 -141
rect -1183 -181 -1171 -147
rect -1133 -181 -1121 -147
rect -1183 -187 -1121 -181
rect -1055 -147 -993 -141
rect -1055 -181 -1043 -147
rect -1005 -181 -993 -147
rect -1055 -187 -993 -181
rect -927 -147 -865 -141
rect -927 -181 -915 -147
rect -877 -181 -865 -147
rect -927 -187 -865 -181
rect -799 -147 -737 -141
rect -799 -181 -787 -147
rect -749 -181 -737 -147
rect -799 -187 -737 -181
rect -671 -147 -609 -141
rect -671 -181 -659 -147
rect -621 -181 -609 -147
rect -671 -187 -609 -181
rect -543 -147 -481 -141
rect -543 -181 -531 -147
rect -493 -181 -481 -147
rect -543 -187 -481 -181
rect -415 -147 -353 -141
rect -415 -181 -403 -147
rect -365 -181 -353 -147
rect -415 -187 -353 -181
rect -287 -147 -225 -141
rect -287 -181 -275 -147
rect -237 -181 -225 -147
rect -287 -187 -225 -181
rect -159 -147 -97 -141
rect -159 -181 -147 -147
rect -109 -181 -97 -147
rect -159 -187 -97 -181
rect -31 -147 31 -141
rect -31 -181 -19 -147
rect 19 -181 31 -147
rect -31 -187 31 -181
rect 97 -147 159 -141
rect 97 -181 109 -147
rect 147 -181 159 -147
rect 97 -187 159 -181
rect 225 -147 287 -141
rect 225 -181 237 -147
rect 275 -181 287 -147
rect 225 -187 287 -181
rect 353 -147 415 -141
rect 353 -181 365 -147
rect 403 -181 415 -147
rect 353 -187 415 -181
rect 481 -147 543 -141
rect 481 -181 493 -147
rect 531 -181 543 -147
rect 481 -187 543 -181
rect 609 -147 671 -141
rect 609 -181 621 -147
rect 659 -181 671 -147
rect 609 -187 671 -181
rect 737 -147 799 -141
rect 737 -181 749 -147
rect 787 -181 799 -147
rect 737 -187 799 -181
rect 865 -147 927 -141
rect 865 -181 877 -147
rect 915 -181 927 -147
rect 865 -187 927 -181
rect 993 -147 1055 -141
rect 993 -181 1005 -147
rect 1043 -181 1055 -147
rect 993 -187 1055 -181
rect 1121 -147 1183 -141
rect 1121 -181 1133 -147
rect 1171 -181 1183 -147
rect 1121 -187 1183 -181
rect 1249 -147 1311 -141
rect 1249 -181 1261 -147
rect 1299 -181 1311 -147
rect 1249 -187 1311 -181
rect 1377 -147 1439 -141
rect 1377 -181 1389 -147
rect 1427 -181 1439 -147
rect 1377 -187 1439 -181
rect 1505 -147 1567 -141
rect 1505 -181 1517 -147
rect 1555 -181 1567 -147
rect 1505 -187 1567 -181
rect 1633 -147 1695 -141
rect 1633 -181 1645 -147
rect 1683 -181 1695 -147
rect 1633 -187 1695 -181
rect 1761 -147 1823 -141
rect 1761 -181 1773 -147
rect 1811 -181 1823 -147
rect 1761 -187 1823 -181
rect 1889 -147 1951 -141
rect 1889 -181 1901 -147
rect 1939 -181 1951 -147
rect 1889 -187 1951 -181
rect 2017 -147 2079 -141
rect 2017 -181 2029 -147
rect 2067 -181 2079 -147
rect 2017 -187 2079 -181
rect 2145 -147 2207 -141
rect 2145 -181 2157 -147
rect 2195 -181 2207 -147
rect 2145 -187 2207 -181
rect 2273 -147 2335 -141
rect 2273 -181 2285 -147
rect 2323 -181 2335 -147
rect 2273 -187 2335 -181
rect 2401 -147 2463 -141
rect 2401 -181 2413 -147
rect 2451 -181 2463 -147
rect 2401 -187 2463 -181
rect 2529 -147 2591 -141
rect 2529 -181 2541 -147
rect 2579 -181 2591 -147
rect 2529 -187 2591 -181
rect 2657 -147 2719 -141
rect 2657 -181 2669 -147
rect 2707 -181 2719 -147
rect 2657 -187 2719 -181
rect 2785 -147 2847 -141
rect 2785 -181 2797 -147
rect 2835 -181 2847 -147
rect 2785 -187 2847 -181
<< properties >>
string FIXED_BBOX -2994 -266 2994 266
string gencell sky130_fd_pr__pfet_01v8_lvt
string library sky130
string parameters w 1.0 l 0.35 m 1 nf 45 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.35 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
