magic
tech sky130A
magscale 1 2
timestamp 1671746218
<< metal3 >>
rect -1350 -900 1349 900
<< mimcap >>
rect -1250 760 1150 800
rect -1250 -760 -1210 760
rect 1110 -760 1150 760
rect -1250 -800 1150 -760
<< mimcapcontact >>
rect -1210 -760 1110 760
<< metal4 >>
rect -1211 760 1111 761
rect -1211 -760 -1210 760
rect 1110 -760 1111 760
rect -1211 -761 1111 -760
<< properties >>
string FIXED_BBOX -1350 -900 1250 900
string gencell sky130_fd_pr__cap_mim_m3_1
string library sky130
string parameters w 12.0 l 8.0 val 199.6 carea 2.00 cperi 0.19 nx 1 ny 1 dummy 0 square 0 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 1 tconnect 1 ccov 100
<< end >>
