magic
tech sky130A
magscale 1 2
timestamp 1672344016
<< nwell >>
rect -957 -1866 957 1866
<< pmoslvt >>
rect -761 118 -661 1718
rect -603 118 -503 1718
rect -445 118 -345 1718
rect -287 118 -187 1718
rect -129 118 -29 1718
rect 29 118 129 1718
rect 187 118 287 1718
rect 345 118 445 1718
rect 503 118 603 1718
rect 661 118 761 1718
rect -761 -1647 -661 -47
rect -603 -1647 -503 -47
rect -445 -1647 -345 -47
rect -287 -1647 -187 -47
rect -129 -1647 -29 -47
rect 29 -1647 129 -47
rect 187 -1647 287 -47
rect 345 -1647 445 -47
rect 503 -1647 603 -47
rect 661 -1647 761 -47
<< pdiff >>
rect -819 1706 -761 1718
rect -819 130 -807 1706
rect -773 130 -761 1706
rect -819 118 -761 130
rect -661 1706 -603 1718
rect -661 130 -649 1706
rect -615 130 -603 1706
rect -661 118 -603 130
rect -503 1706 -445 1718
rect -503 130 -491 1706
rect -457 130 -445 1706
rect -503 118 -445 130
rect -345 1706 -287 1718
rect -345 130 -333 1706
rect -299 130 -287 1706
rect -345 118 -287 130
rect -187 1706 -129 1718
rect -187 130 -175 1706
rect -141 130 -129 1706
rect -187 118 -129 130
rect -29 1706 29 1718
rect -29 130 -17 1706
rect 17 130 29 1706
rect -29 118 29 130
rect 129 1706 187 1718
rect 129 130 141 1706
rect 175 130 187 1706
rect 129 118 187 130
rect 287 1706 345 1718
rect 287 130 299 1706
rect 333 130 345 1706
rect 287 118 345 130
rect 445 1706 503 1718
rect 445 130 457 1706
rect 491 130 503 1706
rect 445 118 503 130
rect 603 1706 661 1718
rect 603 130 615 1706
rect 649 130 661 1706
rect 603 118 661 130
rect 761 1706 819 1718
rect 761 130 773 1706
rect 807 130 819 1706
rect 761 118 819 130
rect -819 -59 -761 -47
rect -819 -1635 -807 -59
rect -773 -1635 -761 -59
rect -819 -1647 -761 -1635
rect -661 -59 -603 -47
rect -661 -1635 -649 -59
rect -615 -1635 -603 -59
rect -661 -1647 -603 -1635
rect -503 -59 -445 -47
rect -503 -1635 -491 -59
rect -457 -1635 -445 -59
rect -503 -1647 -445 -1635
rect -345 -59 -287 -47
rect -345 -1635 -333 -59
rect -299 -1635 -287 -59
rect -345 -1647 -287 -1635
rect -187 -59 -129 -47
rect -187 -1635 -175 -59
rect -141 -1635 -129 -59
rect -187 -1647 -129 -1635
rect -29 -59 29 -47
rect -29 -1635 -17 -59
rect 17 -1635 29 -59
rect -29 -1647 29 -1635
rect 129 -59 187 -47
rect 129 -1635 141 -59
rect 175 -1635 187 -59
rect 129 -1647 187 -1635
rect 287 -59 345 -47
rect 287 -1635 299 -59
rect 333 -1635 345 -59
rect 287 -1647 345 -1635
rect 445 -59 503 -47
rect 445 -1635 457 -59
rect 491 -1635 503 -59
rect 445 -1647 503 -1635
rect 603 -59 661 -47
rect 603 -1635 615 -59
rect 649 -1635 661 -59
rect 603 -1647 661 -1635
rect 761 -59 819 -47
rect 761 -1635 773 -59
rect 807 -1635 819 -59
rect 761 -1647 819 -1635
<< pdiffc >>
rect -807 130 -773 1706
rect -649 130 -615 1706
rect -491 130 -457 1706
rect -333 130 -299 1706
rect -175 130 -141 1706
rect -17 130 17 1706
rect 141 130 175 1706
rect 299 130 333 1706
rect 457 130 491 1706
rect 615 130 649 1706
rect 773 130 807 1706
rect -807 -1635 -773 -59
rect -649 -1635 -615 -59
rect -491 -1635 -457 -59
rect -333 -1635 -299 -59
rect -175 -1635 -141 -59
rect -17 -1635 17 -59
rect 141 -1635 175 -59
rect 299 -1635 333 -59
rect 457 -1635 491 -59
rect 615 -1635 649 -59
rect 773 -1635 807 -59
<< nsubdiff >>
rect -921 1796 -825 1830
rect 825 1796 921 1830
rect -921 1734 -887 1796
rect 887 1734 921 1796
rect -921 -1796 -887 -1734
rect 887 -1796 921 -1734
rect -921 -1830 -825 -1796
rect 825 -1830 921 -1796
<< nsubdiffcont >>
rect -825 1796 825 1830
rect -921 -1734 -887 1734
rect 887 -1734 921 1734
rect -825 -1830 825 -1796
<< poly >>
rect -761 1718 -661 1744
rect -603 1718 -503 1744
rect -445 1718 -345 1744
rect -287 1718 -187 1744
rect -129 1718 -29 1744
rect 29 1718 129 1744
rect 187 1718 287 1744
rect 345 1718 445 1744
rect 503 1718 603 1744
rect 661 1718 761 1744
rect -761 71 -661 118
rect -761 37 -745 71
rect -677 37 -661 71
rect -761 21 -661 37
rect -603 71 -503 118
rect -603 37 -587 71
rect -519 37 -503 71
rect -603 21 -503 37
rect -445 71 -345 118
rect -445 37 -429 71
rect -361 37 -345 71
rect -445 21 -345 37
rect -287 71 -187 118
rect -287 37 -271 71
rect -203 37 -187 71
rect -287 21 -187 37
rect -129 71 -29 118
rect -129 37 -113 71
rect -45 37 -29 71
rect -129 21 -29 37
rect 29 71 129 118
rect 29 37 45 71
rect 113 37 129 71
rect 29 21 129 37
rect 187 71 287 118
rect 187 37 203 71
rect 271 37 287 71
rect 187 21 287 37
rect 345 71 445 118
rect 345 37 361 71
rect 429 37 445 71
rect 345 21 445 37
rect 503 71 603 118
rect 503 37 519 71
rect 587 37 603 71
rect 503 21 603 37
rect 661 71 761 118
rect 661 37 677 71
rect 745 37 761 71
rect 661 21 761 37
rect -761 -47 -661 -21
rect -603 -47 -503 -21
rect -445 -47 -345 -21
rect -287 -47 -187 -21
rect -129 -47 -29 -21
rect 29 -47 129 -21
rect 187 -47 287 -21
rect 345 -47 445 -21
rect 503 -47 603 -21
rect 661 -47 761 -21
rect -761 -1694 -661 -1647
rect -761 -1728 -745 -1694
rect -677 -1728 -661 -1694
rect -761 -1744 -661 -1728
rect -603 -1694 -503 -1647
rect -603 -1728 -587 -1694
rect -519 -1728 -503 -1694
rect -603 -1744 -503 -1728
rect -445 -1694 -345 -1647
rect -445 -1728 -429 -1694
rect -361 -1728 -345 -1694
rect -445 -1744 -345 -1728
rect -287 -1694 -187 -1647
rect -287 -1728 -271 -1694
rect -203 -1728 -187 -1694
rect -287 -1744 -187 -1728
rect -129 -1694 -29 -1647
rect -129 -1728 -113 -1694
rect -45 -1728 -29 -1694
rect -129 -1744 -29 -1728
rect 29 -1694 129 -1647
rect 29 -1728 45 -1694
rect 113 -1728 129 -1694
rect 29 -1744 129 -1728
rect 187 -1694 287 -1647
rect 187 -1728 203 -1694
rect 271 -1728 287 -1694
rect 187 -1744 287 -1728
rect 345 -1694 445 -1647
rect 345 -1728 361 -1694
rect 429 -1728 445 -1694
rect 345 -1744 445 -1728
rect 503 -1694 603 -1647
rect 503 -1728 519 -1694
rect 587 -1728 603 -1694
rect 503 -1744 603 -1728
rect 661 -1694 761 -1647
rect 661 -1728 677 -1694
rect 745 -1728 761 -1694
rect 661 -1744 761 -1728
<< polycont >>
rect -745 37 -677 71
rect -587 37 -519 71
rect -429 37 -361 71
rect -271 37 -203 71
rect -113 37 -45 71
rect 45 37 113 71
rect 203 37 271 71
rect 361 37 429 71
rect 519 37 587 71
rect 677 37 745 71
rect -745 -1728 -677 -1694
rect -587 -1728 -519 -1694
rect -429 -1728 -361 -1694
rect -271 -1728 -203 -1694
rect -113 -1728 -45 -1694
rect 45 -1728 113 -1694
rect 203 -1728 271 -1694
rect 361 -1728 429 -1694
rect 519 -1728 587 -1694
rect 677 -1728 745 -1694
<< locali >>
rect -921 1796 -825 1830
rect 825 1796 921 1830
rect -921 1734 -887 1796
rect 887 1734 921 1796
rect -807 1706 -773 1722
rect -807 114 -773 130
rect -649 1706 -615 1722
rect -649 114 -615 130
rect -491 1706 -457 1722
rect -491 114 -457 130
rect -333 1706 -299 1722
rect -333 114 -299 130
rect -175 1706 -141 1722
rect -175 114 -141 130
rect -17 1706 17 1722
rect -17 114 17 130
rect 141 1706 175 1722
rect 141 114 175 130
rect 299 1706 333 1722
rect 299 114 333 130
rect 457 1706 491 1722
rect 457 114 491 130
rect 615 1706 649 1722
rect 615 114 649 130
rect 773 1706 807 1722
rect 773 114 807 130
rect -761 37 -745 71
rect -677 37 -661 71
rect -603 37 -587 71
rect -519 37 -503 71
rect -445 37 -429 71
rect -361 37 -345 71
rect -287 37 -271 71
rect -203 37 -187 71
rect -129 37 -113 71
rect -45 37 -29 71
rect 29 37 45 71
rect 113 37 129 71
rect 187 37 203 71
rect 271 37 287 71
rect 345 37 361 71
rect 429 37 445 71
rect 503 37 519 71
rect 587 37 603 71
rect 661 37 677 71
rect 745 37 761 71
rect -807 -59 -773 -43
rect -807 -1651 -773 -1635
rect -649 -59 -615 -43
rect -649 -1651 -615 -1635
rect -491 -59 -457 -43
rect -491 -1651 -457 -1635
rect -333 -59 -299 -43
rect -333 -1651 -299 -1635
rect -175 -59 -141 -43
rect -175 -1651 -141 -1635
rect -17 -59 17 -43
rect -17 -1651 17 -1635
rect 141 -59 175 -43
rect 141 -1651 175 -1635
rect 299 -59 333 -43
rect 299 -1651 333 -1635
rect 457 -59 491 -43
rect 457 -1651 491 -1635
rect 615 -59 649 -43
rect 615 -1651 649 -1635
rect 773 -59 807 -43
rect 773 -1651 807 -1635
rect -761 -1728 -745 -1694
rect -677 -1728 -661 -1694
rect -603 -1728 -587 -1694
rect -519 -1728 -503 -1694
rect -445 -1728 -429 -1694
rect -361 -1728 -345 -1694
rect -287 -1728 -271 -1694
rect -203 -1728 -187 -1694
rect -129 -1728 -113 -1694
rect -45 -1728 -29 -1694
rect 29 -1728 45 -1694
rect 113 -1728 129 -1694
rect 187 -1728 203 -1694
rect 271 -1728 287 -1694
rect 345 -1728 361 -1694
rect 429 -1728 445 -1694
rect 503 -1728 519 -1694
rect 587 -1728 603 -1694
rect 661 -1728 677 -1694
rect 745 -1728 761 -1694
rect -921 -1796 -887 -1734
rect 887 -1796 921 -1734
rect -921 -1830 -825 -1796
rect 825 -1830 921 -1796
<< viali >>
rect -807 130 -773 1706
rect -649 130 -615 1706
rect -491 130 -457 1706
rect -333 130 -299 1706
rect -175 130 -141 1706
rect -17 130 17 1706
rect 141 130 175 1706
rect 299 130 333 1706
rect 457 130 491 1706
rect 615 130 649 1706
rect 773 130 807 1706
rect -745 37 -677 71
rect -587 37 -519 71
rect -429 37 -361 71
rect -271 37 -203 71
rect -113 37 -45 71
rect 45 37 113 71
rect 203 37 271 71
rect 361 37 429 71
rect 519 37 587 71
rect 677 37 745 71
rect -807 -1635 -773 -59
rect -649 -1635 -615 -59
rect -491 -1635 -457 -59
rect -333 -1635 -299 -59
rect -175 -1635 -141 -59
rect -17 -1635 17 -59
rect 141 -1635 175 -59
rect 299 -1635 333 -59
rect 457 -1635 491 -59
rect 615 -1635 649 -59
rect 773 -1635 807 -59
rect -745 -1728 -677 -1694
rect -587 -1728 -519 -1694
rect -429 -1728 -361 -1694
rect -271 -1728 -203 -1694
rect -113 -1728 -45 -1694
rect 45 -1728 113 -1694
rect 203 -1728 271 -1694
rect 361 -1728 429 -1694
rect 519 -1728 587 -1694
rect 677 -1728 745 -1694
<< metal1 >>
rect -813 1706 -767 1718
rect -813 130 -807 1706
rect -773 130 -767 1706
rect -813 118 -767 130
rect -655 1706 -609 1718
rect -655 130 -649 1706
rect -615 130 -609 1706
rect -655 118 -609 130
rect -497 1706 -451 1718
rect -497 130 -491 1706
rect -457 130 -451 1706
rect -497 118 -451 130
rect -339 1706 -293 1718
rect -339 130 -333 1706
rect -299 130 -293 1706
rect -339 118 -293 130
rect -181 1706 -135 1718
rect -181 130 -175 1706
rect -141 130 -135 1706
rect -181 118 -135 130
rect -23 1706 23 1718
rect -23 130 -17 1706
rect 17 130 23 1706
rect -23 118 23 130
rect 135 1706 181 1718
rect 135 130 141 1706
rect 175 130 181 1706
rect 135 118 181 130
rect 293 1706 339 1718
rect 293 130 299 1706
rect 333 130 339 1706
rect 293 118 339 130
rect 451 1706 497 1718
rect 451 130 457 1706
rect 491 130 497 1706
rect 451 118 497 130
rect 609 1706 655 1718
rect 609 130 615 1706
rect 649 130 655 1706
rect 609 118 655 130
rect 767 1706 813 1718
rect 767 130 773 1706
rect 807 130 813 1706
rect 767 118 813 130
rect -757 71 -665 77
rect -757 37 -745 71
rect -677 37 -665 71
rect -757 31 -665 37
rect -599 71 -507 77
rect -599 37 -587 71
rect -519 37 -507 71
rect -599 31 -507 37
rect -441 71 -349 77
rect -441 37 -429 71
rect -361 37 -349 71
rect -441 31 -349 37
rect -283 71 -191 77
rect -283 37 -271 71
rect -203 37 -191 71
rect -283 31 -191 37
rect -125 71 -33 77
rect -125 37 -113 71
rect -45 37 -33 71
rect -125 31 -33 37
rect 33 71 125 77
rect 33 37 45 71
rect 113 37 125 71
rect 33 31 125 37
rect 191 71 283 77
rect 191 37 203 71
rect 271 37 283 71
rect 191 31 283 37
rect 349 71 441 77
rect 349 37 361 71
rect 429 37 441 71
rect 349 31 441 37
rect 507 71 599 77
rect 507 37 519 71
rect 587 37 599 71
rect 507 31 599 37
rect 665 71 757 77
rect 665 37 677 71
rect 745 37 757 71
rect 665 31 757 37
rect -813 -59 -767 -47
rect -813 -1635 -807 -59
rect -773 -1635 -767 -59
rect -813 -1647 -767 -1635
rect -655 -59 -609 -47
rect -655 -1635 -649 -59
rect -615 -1635 -609 -59
rect -655 -1647 -609 -1635
rect -497 -59 -451 -47
rect -497 -1635 -491 -59
rect -457 -1635 -451 -59
rect -497 -1647 -451 -1635
rect -339 -59 -293 -47
rect -339 -1635 -333 -59
rect -299 -1635 -293 -59
rect -339 -1647 -293 -1635
rect -181 -59 -135 -47
rect -181 -1635 -175 -59
rect -141 -1635 -135 -59
rect -181 -1647 -135 -1635
rect -23 -59 23 -47
rect -23 -1635 -17 -59
rect 17 -1635 23 -59
rect -23 -1647 23 -1635
rect 135 -59 181 -47
rect 135 -1635 141 -59
rect 175 -1635 181 -59
rect 135 -1647 181 -1635
rect 293 -59 339 -47
rect 293 -1635 299 -59
rect 333 -1635 339 -59
rect 293 -1647 339 -1635
rect 451 -59 497 -47
rect 451 -1635 457 -59
rect 491 -1635 497 -59
rect 451 -1647 497 -1635
rect 609 -59 655 -47
rect 609 -1635 615 -59
rect 649 -1635 655 -59
rect 609 -1647 655 -1635
rect 767 -59 813 -47
rect 767 -1635 773 -59
rect 807 -1635 813 -59
rect 767 -1647 813 -1635
rect -757 -1694 -665 -1688
rect -757 -1728 -745 -1694
rect -677 -1728 -665 -1694
rect -757 -1734 -665 -1728
rect -599 -1694 -507 -1688
rect -599 -1728 -587 -1694
rect -519 -1728 -507 -1694
rect -599 -1734 -507 -1728
rect -441 -1694 -349 -1688
rect -441 -1728 -429 -1694
rect -361 -1728 -349 -1694
rect -441 -1734 -349 -1728
rect -283 -1694 -191 -1688
rect -283 -1728 -271 -1694
rect -203 -1728 -191 -1694
rect -283 -1734 -191 -1728
rect -125 -1694 -33 -1688
rect -125 -1728 -113 -1694
rect -45 -1728 -33 -1694
rect -125 -1734 -33 -1728
rect 33 -1694 125 -1688
rect 33 -1728 45 -1694
rect 113 -1728 125 -1694
rect 33 -1734 125 -1728
rect 191 -1694 283 -1688
rect 191 -1728 203 -1694
rect 271 -1728 283 -1694
rect 191 -1734 283 -1728
rect 349 -1694 441 -1688
rect 349 -1728 361 -1694
rect 429 -1728 441 -1694
rect 349 -1734 441 -1728
rect 507 -1694 599 -1688
rect 507 -1728 519 -1694
rect 587 -1728 599 -1694
rect 507 -1734 599 -1728
rect 665 -1694 757 -1688
rect 665 -1728 677 -1694
rect 745 -1728 757 -1694
rect 665 -1734 757 -1728
<< properties >>
string FIXED_BBOX -904 -1813 904 1813
string gencell sky130_fd_pr__pfet_01v8_lvt
string library sky130
string parameters w 8 l 0.5 m 2 nf 10 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 0 botc 1 poverlap 0 doverlap 1 lmin 0.35 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
