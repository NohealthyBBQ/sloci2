magic
tech sky130A
magscale 1 2
timestamp 1662675866
<< nwell >>
rect -700 -500 2900 3100
<< nsubdiff >>
rect -500 2900 800 3000
rect 1500 2900 2700 3000
rect -500 1700 -400 2900
rect -500 -300 -400 900
rect 2600 1700 2700 2900
rect 2600 -300 2700 900
rect -500 -400 800 -300
rect 1500 -400 2700 -300
<< nsubdiffcont >>
rect 800 2900 1500 3000
rect -500 900 -400 1700
rect 2600 900 2700 1700
rect 800 -400 1500 -300
<< locali >>
rect -500 2900 800 3000
rect 1500 2900 2700 3000
rect -500 1700 -400 2900
rect -500 -300 -400 900
rect 2600 1700 2700 2900
rect 2600 -300 2700 900
rect -500 -400 800 -300
rect 1500 -400 2700 -300
<< metal1 >>
rect 790 2440 800 2500
rect 860 2440 870 2500
rect 1830 2440 1840 2500
rect 1900 2440 1910 2500
rect 30 2360 40 2420
rect 100 2360 110 2420
rect 550 2360 560 2420
rect 620 2360 630 2420
rect 1050 2360 1060 2420
rect 1120 2360 1130 2420
rect 1570 2360 1580 2420
rect 1640 2360 1650 2420
rect 2090 2360 2100 2420
rect 2160 2360 2170 2420
rect 290 2300 300 2360
rect 360 2300 370 2360
rect 1310 2300 1320 2360
rect 1380 2300 1390 2360
rect 98 2202 2096 2250
rect 790 2060 800 2120
rect 860 2060 870 2120
rect 1830 2060 1840 2120
rect 1900 2060 1910 2120
rect 30 2000 40 2060
rect 100 2000 110 2060
rect 550 2000 560 2060
rect 620 2000 630 2060
rect 1050 2000 1060 2060
rect 1120 2000 1130 2060
rect 1570 2000 1580 2060
rect 1640 2000 1650 2060
rect 290 1920 300 1980
rect 360 1920 370 1980
rect 1310 1920 1320 1980
rect 1380 1920 1390 1980
rect 1980 1884 2020 2202
rect 2090 2000 2100 2060
rect 2160 2000 2170 2060
rect 98 1838 2096 1884
rect 790 1700 800 1760
rect 860 1700 870 1760
rect 1830 1700 1840 1760
rect 1900 1700 1910 1760
rect 30 1640 40 1700
rect 100 1640 110 1700
rect 550 1640 560 1700
rect 620 1640 630 1700
rect 1050 1640 1060 1700
rect 1120 1640 1130 1700
rect 1570 1640 1580 1700
rect 1640 1640 1650 1700
rect 290 1560 300 1620
rect 360 1560 370 1620
rect 1310 1560 1320 1620
rect 1380 1560 1390 1620
rect 1980 1520 2020 1838
rect 2090 1640 2100 1700
rect 2160 1640 2170 1700
rect 98 1472 2096 1520
rect 810 1340 820 1400
rect 880 1340 890 1400
rect 1830 1340 1840 1400
rect 1900 1340 1910 1400
rect 30 1280 40 1340
rect 100 1280 110 1340
rect 550 1280 560 1340
rect 620 1280 630 1340
rect 1050 1280 1060 1340
rect 1120 1280 1130 1340
rect 1570 1280 1580 1340
rect 1640 1280 1650 1340
rect 290 1200 300 1260
rect 360 1200 370 1260
rect 1330 1200 1340 1260
rect 1400 1200 1410 1260
rect 1980 1154 2020 1472
rect 2090 1280 2100 1340
rect 2160 1280 2170 1340
rect 98 1108 2096 1154
rect 790 980 800 1040
rect 860 980 870 1040
rect 1830 980 1840 1040
rect 1900 980 1910 1040
rect 30 900 40 960
rect 100 900 110 960
rect 550 900 560 960
rect 620 900 630 960
rect 1050 900 1060 960
rect 1120 900 1130 960
rect 1570 900 1580 960
rect 1640 900 1650 960
rect 290 840 300 900
rect 360 840 370 900
rect 1310 840 1320 900
rect 1380 840 1390 900
rect 1980 790 2020 1108
rect 2090 900 2100 960
rect 2160 900 2170 960
rect 98 742 2096 790
rect 790 600 800 660
rect 860 600 870 660
rect 1830 600 1840 660
rect 1900 600 1910 660
rect 30 540 40 600
rect 100 540 110 600
rect 550 540 560 600
rect 620 540 630 600
rect 1050 540 1060 600
rect 1120 540 1130 600
rect 1570 540 1580 600
rect 1640 540 1650 600
rect 290 460 300 520
rect 360 460 370 520
rect 1310 460 1320 520
rect 1380 460 1390 520
rect 1980 424 2020 742
rect 2090 540 2100 600
rect 2160 540 2170 600
rect 98 378 2096 424
rect 790 240 800 300
rect 860 240 870 300
rect 1830 240 1840 300
rect 1900 240 1910 300
rect 30 180 40 240
rect 100 180 110 240
rect 550 180 560 240
rect 620 180 630 240
rect 1050 180 1060 240
rect 1120 180 1130 240
rect 1570 180 1580 240
rect 1640 180 1650 240
rect 290 100 300 160
rect 360 100 370 160
rect 1310 100 1320 160
rect 1380 100 1390 160
rect 1980 60 2020 378
rect 2090 180 2100 240
rect 2160 180 2170 240
rect 98 12 2096 60
<< via1 >>
rect 800 2440 860 2500
rect 1840 2440 1900 2500
rect 40 2360 100 2420
rect 560 2360 620 2420
rect 1060 2360 1120 2420
rect 1580 2360 1640 2420
rect 2100 2360 2160 2420
rect 300 2300 360 2360
rect 1320 2300 1380 2360
rect 800 2060 860 2120
rect 1840 2060 1900 2120
rect 40 2000 100 2060
rect 560 2000 620 2060
rect 1060 2000 1120 2060
rect 1580 2000 1640 2060
rect 300 1920 360 1980
rect 1320 1920 1380 1980
rect 2100 2000 2160 2060
rect 800 1700 860 1760
rect 1840 1700 1900 1760
rect 40 1640 100 1700
rect 560 1640 620 1700
rect 1060 1640 1120 1700
rect 1580 1640 1640 1700
rect 300 1560 360 1620
rect 1320 1560 1380 1620
rect 2100 1640 2160 1700
rect 820 1340 880 1400
rect 1840 1340 1900 1400
rect 40 1280 100 1340
rect 560 1280 620 1340
rect 1060 1280 1120 1340
rect 1580 1280 1640 1340
rect 300 1200 360 1260
rect 1340 1200 1400 1260
rect 2100 1280 2160 1340
rect 800 980 860 1040
rect 1840 980 1900 1040
rect 40 900 100 960
rect 560 900 620 960
rect 1060 900 1120 960
rect 1580 900 1640 960
rect 300 840 360 900
rect 1320 840 1380 900
rect 2100 900 2160 960
rect 800 600 860 660
rect 1840 600 1900 660
rect 40 540 100 600
rect 560 540 620 600
rect 1060 540 1120 600
rect 1580 540 1640 600
rect 300 460 360 520
rect 1320 460 1380 520
rect 2100 540 2160 600
rect 800 240 860 300
rect 1840 240 1900 300
rect 40 180 100 240
rect 560 180 620 240
rect 1060 180 1120 240
rect 1580 180 1640 240
rect 300 100 360 160
rect 1320 100 1380 160
rect 2100 180 2160 240
<< metal2 >>
rect 800 2500 2320 2520
rect 860 2480 1840 2500
rect 800 2430 860 2440
rect 1900 2480 2320 2500
rect 1840 2430 1900 2440
rect 40 2420 100 2430
rect 560 2420 620 2430
rect 40 2350 100 2360
rect 300 2360 360 2370
rect -120 2300 300 2320
rect 560 2350 620 2360
rect 1060 2420 1120 2430
rect 1580 2420 1640 2430
rect 1060 2350 1120 2360
rect 1320 2360 1380 2370
rect 360 2300 1320 2320
rect 1580 2350 1640 2360
rect 2100 2420 2160 2430
rect 2100 2350 2160 2360
rect -120 2280 1380 2300
rect -120 2140 -40 2280
rect -120 2120 1900 2140
rect -120 2100 800 2120
rect -120 1580 -40 2100
rect 40 2060 100 2070
rect 40 1990 100 2000
rect 560 2060 620 2070
rect 860 2100 1840 2120
rect 800 2050 860 2060
rect 1060 2060 1120 2070
rect 560 1990 620 2000
rect 1060 1990 1120 2000
rect 1580 2060 1640 2070
rect 1840 2050 1900 2060
rect 2100 2060 2160 2070
rect 1580 1990 1640 2000
rect 2100 1990 2160 2000
rect 300 1980 360 1990
rect 1320 1980 1380 1990
rect 360 1920 1320 1940
rect 2240 1940 2320 2480
rect 1380 1920 2320 1940
rect 300 1900 2320 1920
rect 2240 1780 2320 1900
rect 800 1760 2320 1780
rect 40 1700 100 1710
rect 40 1630 100 1640
rect 560 1700 620 1710
rect 860 1740 1840 1760
rect 800 1690 860 1700
rect 1060 1700 1120 1710
rect 560 1630 620 1640
rect 1060 1630 1120 1640
rect 1580 1700 1640 1710
rect 1900 1740 2320 1760
rect 1840 1690 1900 1700
rect 2100 1700 2160 1710
rect 1580 1630 1640 1640
rect 2100 1630 2160 1640
rect 300 1620 360 1630
rect -120 1560 300 1580
rect 1320 1620 1380 1630
rect 360 1560 1320 1580
rect -120 1540 1380 1560
rect -120 1420 -40 1540
rect -120 1400 1900 1420
rect -120 1380 820 1400
rect -120 860 -40 1380
rect 40 1340 100 1350
rect 40 1270 100 1280
rect 560 1340 620 1350
rect 880 1380 1840 1400
rect 820 1330 880 1340
rect 1060 1340 1120 1350
rect 560 1270 620 1280
rect 1060 1270 1120 1280
rect 1580 1340 1640 1350
rect 1840 1330 1900 1340
rect 2100 1340 2160 1350
rect 1580 1270 1640 1280
rect 2100 1270 2160 1280
rect 300 1260 360 1270
rect 1340 1260 1400 1270
rect 360 1200 1340 1220
rect 2240 1220 2320 1740
rect 1400 1200 2320 1220
rect 300 1180 2320 1200
rect 2240 1060 2320 1180
rect 800 1040 2320 1060
rect 860 1020 1840 1040
rect 800 970 860 980
rect 1900 1020 2320 1040
rect 1840 970 1900 980
rect 40 960 100 970
rect 560 960 620 970
rect 40 890 100 900
rect 300 900 360 910
rect -120 840 300 860
rect 560 890 620 900
rect 1060 960 1120 970
rect 1580 960 1640 970
rect 1060 890 1120 900
rect 1320 900 1380 910
rect 360 840 1320 860
rect 1580 890 1640 900
rect 2100 960 2160 970
rect 2100 890 2160 900
rect -120 820 1380 840
rect -120 680 -40 820
rect -120 660 1900 680
rect -120 640 800 660
rect -120 120 -40 640
rect 40 600 100 610
rect 40 530 100 540
rect 560 600 620 610
rect 860 640 1840 660
rect 800 590 860 600
rect 1060 600 1120 610
rect 560 530 620 540
rect 1060 530 1120 540
rect 1580 600 1640 610
rect 1840 590 1900 600
rect 2100 600 2160 610
rect 1580 530 1640 540
rect 2100 530 2160 540
rect 300 520 360 530
rect 1320 520 1380 530
rect 360 460 1320 480
rect 2240 480 2320 1020
rect 1380 460 2320 480
rect 300 440 2320 460
rect 2240 320 2320 440
rect 800 300 2320 320
rect 40 240 100 250
rect 40 170 100 180
rect 560 240 620 250
rect 860 280 1840 300
rect 800 230 860 240
rect 1060 240 1120 250
rect 560 170 620 180
rect 1060 170 1120 180
rect 1580 240 1640 250
rect 1900 280 2320 300
rect 1840 230 1900 240
rect 2100 240 2160 250
rect 1580 170 1640 180
rect 2100 170 2160 180
rect 300 160 360 170
rect -120 100 300 120
rect 1320 160 1380 170
rect 360 100 1320 120
rect -120 80 1380 100
<< via2 >>
rect 40 2360 100 2420
rect 560 2360 620 2420
rect 1060 2360 1120 2420
rect 1580 2360 1640 2420
rect 2100 2360 2160 2420
rect 40 2000 100 2060
rect 560 2000 620 2060
rect 1060 2000 1120 2060
rect 1580 2000 1640 2060
rect 2100 2000 2160 2060
rect 40 1640 100 1700
rect 560 1640 620 1700
rect 1060 1640 1120 1700
rect 1580 1640 1640 1700
rect 2100 1640 2160 1700
rect 40 1280 100 1340
rect 560 1280 620 1340
rect 1060 1280 1120 1340
rect 1580 1280 1640 1340
rect 2100 1280 2160 1340
rect 40 900 100 960
rect 560 900 620 960
rect 1060 900 1120 960
rect 1580 900 1640 960
rect 2100 900 2160 960
rect 40 540 100 600
rect 560 540 620 600
rect 1060 540 1120 600
rect 1580 540 1640 600
rect 2100 540 2160 600
rect 40 180 100 240
rect 560 180 620 240
rect 1060 180 1120 240
rect 1580 180 1640 240
rect 2100 180 2160 240
<< metal3 >>
rect 40 2425 100 2500
rect 560 2425 620 2500
rect 1060 2425 1120 2500
rect 1580 2425 1640 2500
rect 2100 2425 2160 2500
rect 30 2420 110 2425
rect 30 2360 40 2420
rect 100 2360 110 2420
rect 30 2355 110 2360
rect 550 2420 630 2425
rect 550 2360 560 2420
rect 620 2360 630 2420
rect 550 2355 630 2360
rect 1050 2420 1130 2425
rect 1050 2360 1060 2420
rect 1120 2360 1130 2420
rect 1050 2355 1130 2360
rect 1570 2420 1650 2425
rect 1570 2360 1580 2420
rect 1640 2360 1650 2420
rect 1570 2355 1650 2360
rect 2090 2420 2170 2425
rect 2090 2360 2100 2420
rect 2160 2360 2170 2420
rect 2090 2355 2170 2360
rect 40 2065 100 2355
rect 560 2065 620 2355
rect 1060 2065 1120 2355
rect 1580 2065 1640 2355
rect 2100 2065 2160 2355
rect 30 2060 110 2065
rect 30 2000 40 2060
rect 100 2000 110 2060
rect 30 1995 110 2000
rect 550 2060 630 2065
rect 550 2000 560 2060
rect 620 2000 630 2060
rect 550 1995 630 2000
rect 1050 2060 1130 2065
rect 1050 2000 1060 2060
rect 1120 2000 1130 2060
rect 1050 1995 1130 2000
rect 1570 2060 1650 2065
rect 1570 2000 1580 2060
rect 1640 2000 1650 2060
rect 1570 1995 1650 2000
rect 2090 2060 2170 2065
rect 2090 2000 2100 2060
rect 2160 2000 2170 2060
rect 2090 1995 2170 2000
rect 40 1705 100 1995
rect 560 1705 620 1995
rect 1060 1705 1120 1995
rect 1580 1705 1640 1995
rect 2100 1705 2160 1995
rect 30 1700 110 1705
rect 30 1640 40 1700
rect 100 1640 110 1700
rect 30 1635 110 1640
rect 550 1700 630 1705
rect 550 1640 560 1700
rect 620 1640 630 1700
rect 550 1635 630 1640
rect 1050 1700 1130 1705
rect 1050 1640 1060 1700
rect 1120 1640 1130 1700
rect 1050 1635 1130 1640
rect 1570 1700 1650 1705
rect 1570 1640 1580 1700
rect 1640 1640 1650 1700
rect 1570 1635 1650 1640
rect 2090 1700 2170 1705
rect 2090 1640 2100 1700
rect 2160 1640 2170 1700
rect 2090 1635 2170 1640
rect 40 1345 100 1635
rect 560 1345 620 1635
rect 1060 1345 1120 1635
rect 1580 1345 1640 1635
rect 2100 1345 2160 1635
rect 30 1340 110 1345
rect 550 1340 630 1345
rect 1050 1340 1130 1345
rect 1570 1340 1650 1345
rect 2090 1340 2170 1345
rect -120 1280 40 1340
rect 100 1280 560 1340
rect 620 1280 1060 1340
rect 1120 1280 1580 1340
rect 1640 1280 2100 1340
rect 2160 1280 2320 1340
rect 30 1275 110 1280
rect 550 1275 630 1280
rect 1050 1275 1130 1280
rect 1570 1275 1650 1280
rect 2090 1275 2170 1280
rect 40 965 100 1275
rect 560 965 620 1275
rect 1060 965 1120 1275
rect 1580 965 1640 1275
rect 2100 965 2160 1275
rect 30 960 110 965
rect 30 900 40 960
rect 100 900 110 960
rect 30 895 110 900
rect 550 960 630 965
rect 550 900 560 960
rect 620 900 630 960
rect 550 895 630 900
rect 1050 960 1130 965
rect 1050 900 1060 960
rect 1120 900 1130 960
rect 1050 895 1130 900
rect 1570 960 1650 965
rect 1570 900 1580 960
rect 1640 900 1650 960
rect 1570 895 1650 900
rect 2090 960 2170 965
rect 2090 900 2100 960
rect 2160 900 2170 960
rect 2090 895 2170 900
rect 40 605 100 895
rect 560 605 620 895
rect 1060 605 1120 895
rect 1580 605 1640 895
rect 2100 605 2160 895
rect 30 600 110 605
rect 30 540 40 600
rect 100 540 110 600
rect 30 535 110 540
rect 550 600 630 605
rect 550 540 560 600
rect 620 540 630 600
rect 550 535 630 540
rect 1050 600 1130 605
rect 1050 540 1060 600
rect 1120 540 1130 600
rect 1050 535 1130 540
rect 1570 600 1650 605
rect 1570 540 1580 600
rect 1640 540 1650 600
rect 1570 535 1650 540
rect 2090 600 2170 605
rect 2090 540 2100 600
rect 2160 540 2170 600
rect 2090 535 2170 540
rect 40 245 100 535
rect 560 245 620 535
rect 1060 245 1120 535
rect 1580 245 1640 535
rect 2100 245 2160 535
rect 30 240 110 245
rect 30 180 40 240
rect 100 180 110 240
rect 30 175 110 180
rect 550 240 630 245
rect 550 180 560 240
rect 620 180 630 240
rect 550 175 630 180
rect 1050 240 1130 245
rect 1050 180 1060 240
rect 1120 180 1130 240
rect 1050 175 1130 180
rect 1570 240 1650 245
rect 1570 180 1580 240
rect 1640 180 1650 240
rect 1570 175 1650 180
rect 2090 240 2170 245
rect 2090 180 2100 240
rect 2160 180 2170 240
rect 2090 175 2170 180
rect 40 100 100 175
rect 560 100 620 175
rect 1060 100 1120 175
rect 1580 100 1640 175
rect 2100 100 2160 175
use sky130_fd_pr__pfet_01v8_lvt_8URDWJ  sky130_fd_pr__pfet_01v8_lvt_8URDWJ_0
timestamp 1662671833
transform 1 0 1097 0 1 1260
box -1097 -1260 1097 1292
<< labels >>
flabel nwell 300 2540 360 2620 0 FreeSans 800 0 0 0 A
flabel nwell 1340 2540 1400 2620 0 FreeSans 800 0 0 0 A
flabel nwell 820 2160 880 2240 0 FreeSans 800 0 0 0 A
flabel nwell 1840 2140 1900 2220 0 FreeSans 800 0 0 0 A
flabel nwell 280 1780 340 1860 0 FreeSans 800 0 0 0 A
flabel nwell 1340 1800 1400 1880 0 FreeSans 800 0 0 0 A
flabel nwell 820 1400 880 1480 0 FreeSans 800 0 0 0 A
flabel nwell 1840 1400 1900 1480 0 FreeSans 800 0 0 0 A
flabel nwell 300 1040 360 1120 0 FreeSans 800 0 0 0 A
flabel nwell 1340 1060 1400 1140 0 FreeSans 800 0 0 0 A
flabel nwell 780 680 840 760 0 FreeSans 800 0 0 0 A
flabel nwell 1860 680 1920 760 0 FreeSans 800 0 0 0 A
flabel nwell 280 300 340 380 0 FreeSans 800 0 0 0 A
flabel nwell 1320 300 1380 380 0 FreeSans 800 0 0 0 A
flabel nwell 820 2520 880 2600 0 FreeSans 800 0 0 0 B
flabel nwell 1840 2520 1900 2600 0 FreeSans 800 0 0 0 B
flabel nwell 300 2140 360 2220 0 FreeSans 800 0 0 0 B
flabel nwell 1340 2140 1400 2220 0 FreeSans 800 0 0 0 B
flabel nwell 820 1780 880 1860 0 FreeSans 800 0 0 0 B
flabel nwell 1860 1780 1920 1860 0 FreeSans 800 0 0 0 B
flabel nwell 280 1400 340 1480 0 FreeSans 800 0 0 0 B
flabel nwell 1340 1420 1400 1500 0 FreeSans 800 0 0 0 B
flabel nwell 820 1060 880 1140 0 FreeSans 800 0 0 0 B
flabel nwell 1840 1060 1900 1140 0 FreeSans 800 0 0 0 B
flabel nwell 300 700 360 780 0 FreeSans 800 0 0 0 B
flabel nwell 1340 680 1400 760 0 FreeSans 800 0 0 0 B
flabel nwell 820 320 880 400 0 FreeSans 800 0 0 0 B
flabel nwell 1840 320 1900 400 0 FreeSans 800 0 0 0 B
<< end >>
