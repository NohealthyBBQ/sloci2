magic
tech sky130A
magscale 1 2
timestamp 1662827102
<< pwell >>
rect -307 -5348 307 5348
<< psubdiff >>
rect -271 5278 -175 5312
rect 175 5278 271 5312
rect -271 5216 -237 5278
rect 237 5216 271 5278
rect -271 -5278 -237 -5216
rect 237 -5278 271 -5216
rect -271 -5312 -175 -5278
rect 175 -5312 271 -5278
<< psubdiffcont >>
rect -175 5278 175 5312
rect -271 -5216 -237 5216
rect 237 -5216 271 5216
rect -175 -5312 175 -5278
<< xpolycontact >>
rect -141 4750 141 5182
rect -141 -5182 141 -4750
<< ppolyres >>
rect -141 -4750 141 4750
<< locali >>
rect -271 5278 -175 5312
rect 175 5278 271 5312
rect -271 5216 -237 5278
rect 237 5216 271 5278
rect -271 -5278 -237 -5216
rect 237 -5278 271 -5216
rect -271 -5312 -175 -5278
rect 175 -5312 271 -5278
<< viali >>
rect -125 4767 125 5164
rect -125 -5164 125 -4767
<< metal1 >>
rect -131 5164 131 5176
rect -131 4767 -125 5164
rect 125 4767 131 5164
rect -131 4755 131 4767
rect -131 -4767 131 -4755
rect -131 -5164 -125 -4767
rect 125 -5164 131 -4767
rect -131 -5176 131 -5164
<< res1p41 >>
rect -143 -4752 143 4752
<< properties >>
string FIXED_BBOX -254 -5295 254 5295
string gencell sky130_fd_pr__res_high_po_1p41
string library sky130
string parameters w 1.410 l 47.5 m 1 nx 1 wmin 1.410 lmin 0.50 rho 319.8 val 11.049k dummy 0 dw 0.0 term 194.82 sterm 0.0 caplen 0 guard 1 glc 1 grc 1 gtc 1 gbc 1 compatible {sky130_fd_pr__res_high_po_0p35  sky130_fd_pr__res_high_po_0p69 sky130_fd_pr__res_high_po_1p41  sky130_fd_pr__res_high_po_2p85 sky130_fd_pr__res_high_po_5p73} snake 0 full_metal 1 wmax 1.410 n_guard 0 hv_guard 0 vias 1 viagb 0 viagt 0 viagl 0 viagr 0
<< end >>
