magic
tech sky130A
magscale 1 2
timestamp 1662404926
<< error_p >>
rect -1887 181 -1825 187
rect -1759 181 -1697 187
rect -1631 181 -1569 187
rect -1503 181 -1441 187
rect -1375 181 -1313 187
rect -1247 181 -1185 187
rect -1119 181 -1057 187
rect -991 181 -929 187
rect -863 181 -801 187
rect -735 181 -673 187
rect -607 181 -545 187
rect -479 181 -417 187
rect -351 181 -289 187
rect -223 181 -161 187
rect -95 181 -33 187
rect 33 181 95 187
rect 161 181 223 187
rect 289 181 351 187
rect 417 181 479 187
rect 545 181 607 187
rect 673 181 735 187
rect 801 181 863 187
rect 929 181 991 187
rect 1057 181 1119 187
rect 1185 181 1247 187
rect 1313 181 1375 187
rect 1441 181 1503 187
rect 1569 181 1631 187
rect 1697 181 1759 187
rect 1825 181 1887 187
rect -1887 147 -1875 181
rect -1759 147 -1747 181
rect -1631 147 -1619 181
rect -1503 147 -1491 181
rect -1375 147 -1363 181
rect -1247 147 -1235 181
rect -1119 147 -1107 181
rect -991 147 -979 181
rect -863 147 -851 181
rect -735 147 -723 181
rect -607 147 -595 181
rect -479 147 -467 181
rect -351 147 -339 181
rect -223 147 -211 181
rect -95 147 -83 181
rect 33 147 45 181
rect 161 147 173 181
rect 289 147 301 181
rect 417 147 429 181
rect 545 147 557 181
rect 673 147 685 181
rect 801 147 813 181
rect 929 147 941 181
rect 1057 147 1069 181
rect 1185 147 1197 181
rect 1313 147 1325 181
rect 1441 147 1453 181
rect 1569 147 1581 181
rect 1697 147 1709 181
rect 1825 147 1837 181
rect -1887 141 -1825 147
rect -1759 141 -1697 147
rect -1631 141 -1569 147
rect -1503 141 -1441 147
rect -1375 141 -1313 147
rect -1247 141 -1185 147
rect -1119 141 -1057 147
rect -991 141 -929 147
rect -863 141 -801 147
rect -735 141 -673 147
rect -607 141 -545 147
rect -479 141 -417 147
rect -351 141 -289 147
rect -223 141 -161 147
rect -95 141 -33 147
rect 33 141 95 147
rect 161 141 223 147
rect 289 141 351 147
rect 417 141 479 147
rect 545 141 607 147
rect 673 141 735 147
rect 801 141 863 147
rect 929 141 991 147
rect 1057 141 1119 147
rect 1185 141 1247 147
rect 1313 141 1375 147
rect 1441 141 1503 147
rect 1569 141 1631 147
rect 1697 141 1759 147
rect 1825 141 1887 147
rect -1887 -147 -1825 -141
rect -1759 -147 -1697 -141
rect -1631 -147 -1569 -141
rect -1503 -147 -1441 -141
rect -1375 -147 -1313 -141
rect -1247 -147 -1185 -141
rect -1119 -147 -1057 -141
rect -991 -147 -929 -141
rect -863 -147 -801 -141
rect -735 -147 -673 -141
rect -607 -147 -545 -141
rect -479 -147 -417 -141
rect -351 -147 -289 -141
rect -223 -147 -161 -141
rect -95 -147 -33 -141
rect 33 -147 95 -141
rect 161 -147 223 -141
rect 289 -147 351 -141
rect 417 -147 479 -141
rect 545 -147 607 -141
rect 673 -147 735 -141
rect 801 -147 863 -141
rect 929 -147 991 -141
rect 1057 -147 1119 -141
rect 1185 -147 1247 -141
rect 1313 -147 1375 -141
rect 1441 -147 1503 -141
rect 1569 -147 1631 -141
rect 1697 -147 1759 -141
rect 1825 -147 1887 -141
rect -1887 -181 -1875 -147
rect -1759 -181 -1747 -147
rect -1631 -181 -1619 -147
rect -1503 -181 -1491 -147
rect -1375 -181 -1363 -147
rect -1247 -181 -1235 -147
rect -1119 -181 -1107 -147
rect -991 -181 -979 -147
rect -863 -181 -851 -147
rect -735 -181 -723 -147
rect -607 -181 -595 -147
rect -479 -181 -467 -147
rect -351 -181 -339 -147
rect -223 -181 -211 -147
rect -95 -181 -83 -147
rect 33 -181 45 -147
rect 161 -181 173 -147
rect 289 -181 301 -147
rect 417 -181 429 -147
rect 545 -181 557 -147
rect 673 -181 685 -147
rect 801 -181 813 -147
rect 929 -181 941 -147
rect 1057 -181 1069 -147
rect 1185 -181 1197 -147
rect 1313 -181 1325 -147
rect 1441 -181 1453 -147
rect 1569 -181 1581 -147
rect 1697 -181 1709 -147
rect 1825 -181 1837 -147
rect -1887 -187 -1825 -181
rect -1759 -187 -1697 -181
rect -1631 -187 -1569 -181
rect -1503 -187 -1441 -181
rect -1375 -187 -1313 -181
rect -1247 -187 -1185 -181
rect -1119 -187 -1057 -181
rect -991 -187 -929 -181
rect -863 -187 -801 -181
rect -735 -187 -673 -181
rect -607 -187 -545 -181
rect -479 -187 -417 -181
rect -351 -187 -289 -181
rect -223 -187 -161 -181
rect -95 -187 -33 -181
rect 33 -187 95 -181
rect 161 -187 223 -181
rect 289 -187 351 -181
rect 417 -187 479 -181
rect 545 -187 607 -181
rect 673 -187 735 -181
rect 801 -187 863 -181
rect 929 -187 991 -181
rect 1057 -187 1119 -181
rect 1185 -187 1247 -181
rect 1313 -187 1375 -181
rect 1441 -187 1503 -181
rect 1569 -187 1631 -181
rect 1697 -187 1759 -181
rect 1825 -187 1887 -181
<< nwell >>
rect -2087 -319 2087 319
<< pmoslvt >>
rect -1891 -100 -1821 100
rect -1763 -100 -1693 100
rect -1635 -100 -1565 100
rect -1507 -100 -1437 100
rect -1379 -100 -1309 100
rect -1251 -100 -1181 100
rect -1123 -100 -1053 100
rect -995 -100 -925 100
rect -867 -100 -797 100
rect -739 -100 -669 100
rect -611 -100 -541 100
rect -483 -100 -413 100
rect -355 -100 -285 100
rect -227 -100 -157 100
rect -99 -100 -29 100
rect 29 -100 99 100
rect 157 -100 227 100
rect 285 -100 355 100
rect 413 -100 483 100
rect 541 -100 611 100
rect 669 -100 739 100
rect 797 -100 867 100
rect 925 -100 995 100
rect 1053 -100 1123 100
rect 1181 -100 1251 100
rect 1309 -100 1379 100
rect 1437 -100 1507 100
rect 1565 -100 1635 100
rect 1693 -100 1763 100
rect 1821 -100 1891 100
<< pdiff >>
rect -1949 88 -1891 100
rect -1949 -88 -1937 88
rect -1903 -88 -1891 88
rect -1949 -100 -1891 -88
rect -1821 88 -1763 100
rect -1821 -88 -1809 88
rect -1775 -88 -1763 88
rect -1821 -100 -1763 -88
rect -1693 88 -1635 100
rect -1693 -88 -1681 88
rect -1647 -88 -1635 88
rect -1693 -100 -1635 -88
rect -1565 88 -1507 100
rect -1565 -88 -1553 88
rect -1519 -88 -1507 88
rect -1565 -100 -1507 -88
rect -1437 88 -1379 100
rect -1437 -88 -1425 88
rect -1391 -88 -1379 88
rect -1437 -100 -1379 -88
rect -1309 88 -1251 100
rect -1309 -88 -1297 88
rect -1263 -88 -1251 88
rect -1309 -100 -1251 -88
rect -1181 88 -1123 100
rect -1181 -88 -1169 88
rect -1135 -88 -1123 88
rect -1181 -100 -1123 -88
rect -1053 88 -995 100
rect -1053 -88 -1041 88
rect -1007 -88 -995 88
rect -1053 -100 -995 -88
rect -925 88 -867 100
rect -925 -88 -913 88
rect -879 -88 -867 88
rect -925 -100 -867 -88
rect -797 88 -739 100
rect -797 -88 -785 88
rect -751 -88 -739 88
rect -797 -100 -739 -88
rect -669 88 -611 100
rect -669 -88 -657 88
rect -623 -88 -611 88
rect -669 -100 -611 -88
rect -541 88 -483 100
rect -541 -88 -529 88
rect -495 -88 -483 88
rect -541 -100 -483 -88
rect -413 88 -355 100
rect -413 -88 -401 88
rect -367 -88 -355 88
rect -413 -100 -355 -88
rect -285 88 -227 100
rect -285 -88 -273 88
rect -239 -88 -227 88
rect -285 -100 -227 -88
rect -157 88 -99 100
rect -157 -88 -145 88
rect -111 -88 -99 88
rect -157 -100 -99 -88
rect -29 88 29 100
rect -29 -88 -17 88
rect 17 -88 29 88
rect -29 -100 29 -88
rect 99 88 157 100
rect 99 -88 111 88
rect 145 -88 157 88
rect 99 -100 157 -88
rect 227 88 285 100
rect 227 -88 239 88
rect 273 -88 285 88
rect 227 -100 285 -88
rect 355 88 413 100
rect 355 -88 367 88
rect 401 -88 413 88
rect 355 -100 413 -88
rect 483 88 541 100
rect 483 -88 495 88
rect 529 -88 541 88
rect 483 -100 541 -88
rect 611 88 669 100
rect 611 -88 623 88
rect 657 -88 669 88
rect 611 -100 669 -88
rect 739 88 797 100
rect 739 -88 751 88
rect 785 -88 797 88
rect 739 -100 797 -88
rect 867 88 925 100
rect 867 -88 879 88
rect 913 -88 925 88
rect 867 -100 925 -88
rect 995 88 1053 100
rect 995 -88 1007 88
rect 1041 -88 1053 88
rect 995 -100 1053 -88
rect 1123 88 1181 100
rect 1123 -88 1135 88
rect 1169 -88 1181 88
rect 1123 -100 1181 -88
rect 1251 88 1309 100
rect 1251 -88 1263 88
rect 1297 -88 1309 88
rect 1251 -100 1309 -88
rect 1379 88 1437 100
rect 1379 -88 1391 88
rect 1425 -88 1437 88
rect 1379 -100 1437 -88
rect 1507 88 1565 100
rect 1507 -88 1519 88
rect 1553 -88 1565 88
rect 1507 -100 1565 -88
rect 1635 88 1693 100
rect 1635 -88 1647 88
rect 1681 -88 1693 88
rect 1635 -100 1693 -88
rect 1763 88 1821 100
rect 1763 -88 1775 88
rect 1809 -88 1821 88
rect 1763 -100 1821 -88
rect 1891 88 1949 100
rect 1891 -88 1903 88
rect 1937 -88 1949 88
rect 1891 -100 1949 -88
<< pdiffc >>
rect -1937 -88 -1903 88
rect -1809 -88 -1775 88
rect -1681 -88 -1647 88
rect -1553 -88 -1519 88
rect -1425 -88 -1391 88
rect -1297 -88 -1263 88
rect -1169 -88 -1135 88
rect -1041 -88 -1007 88
rect -913 -88 -879 88
rect -785 -88 -751 88
rect -657 -88 -623 88
rect -529 -88 -495 88
rect -401 -88 -367 88
rect -273 -88 -239 88
rect -145 -88 -111 88
rect -17 -88 17 88
rect 111 -88 145 88
rect 239 -88 273 88
rect 367 -88 401 88
rect 495 -88 529 88
rect 623 -88 657 88
rect 751 -88 785 88
rect 879 -88 913 88
rect 1007 -88 1041 88
rect 1135 -88 1169 88
rect 1263 -88 1297 88
rect 1391 -88 1425 88
rect 1519 -88 1553 88
rect 1647 -88 1681 88
rect 1775 -88 1809 88
rect 1903 -88 1937 88
<< nsubdiff >>
rect -2051 249 -1955 283
rect 1955 249 2051 283
rect -2051 187 -2017 249
rect 2017 187 2051 249
rect -2051 -249 -2017 -187
rect 2017 -249 2051 -187
rect -2051 -283 -1955 -249
rect 1955 -283 2051 -249
<< nsubdiffcont >>
rect -1955 249 1955 283
rect -2051 -187 -2017 187
rect 2017 -187 2051 187
rect -1955 -283 1955 -249
<< poly >>
rect -1891 181 -1821 197
rect -1891 147 -1875 181
rect -1837 147 -1821 181
rect -1891 100 -1821 147
rect -1763 181 -1693 197
rect -1763 147 -1747 181
rect -1709 147 -1693 181
rect -1763 100 -1693 147
rect -1635 181 -1565 197
rect -1635 147 -1619 181
rect -1581 147 -1565 181
rect -1635 100 -1565 147
rect -1507 181 -1437 197
rect -1507 147 -1491 181
rect -1453 147 -1437 181
rect -1507 100 -1437 147
rect -1379 181 -1309 197
rect -1379 147 -1363 181
rect -1325 147 -1309 181
rect -1379 100 -1309 147
rect -1251 181 -1181 197
rect -1251 147 -1235 181
rect -1197 147 -1181 181
rect -1251 100 -1181 147
rect -1123 181 -1053 197
rect -1123 147 -1107 181
rect -1069 147 -1053 181
rect -1123 100 -1053 147
rect -995 181 -925 197
rect -995 147 -979 181
rect -941 147 -925 181
rect -995 100 -925 147
rect -867 181 -797 197
rect -867 147 -851 181
rect -813 147 -797 181
rect -867 100 -797 147
rect -739 181 -669 197
rect -739 147 -723 181
rect -685 147 -669 181
rect -739 100 -669 147
rect -611 181 -541 197
rect -611 147 -595 181
rect -557 147 -541 181
rect -611 100 -541 147
rect -483 181 -413 197
rect -483 147 -467 181
rect -429 147 -413 181
rect -483 100 -413 147
rect -355 181 -285 197
rect -355 147 -339 181
rect -301 147 -285 181
rect -355 100 -285 147
rect -227 181 -157 197
rect -227 147 -211 181
rect -173 147 -157 181
rect -227 100 -157 147
rect -99 181 -29 197
rect -99 147 -83 181
rect -45 147 -29 181
rect -99 100 -29 147
rect 29 181 99 197
rect 29 147 45 181
rect 83 147 99 181
rect 29 100 99 147
rect 157 181 227 197
rect 157 147 173 181
rect 211 147 227 181
rect 157 100 227 147
rect 285 181 355 197
rect 285 147 301 181
rect 339 147 355 181
rect 285 100 355 147
rect 413 181 483 197
rect 413 147 429 181
rect 467 147 483 181
rect 413 100 483 147
rect 541 181 611 197
rect 541 147 557 181
rect 595 147 611 181
rect 541 100 611 147
rect 669 181 739 197
rect 669 147 685 181
rect 723 147 739 181
rect 669 100 739 147
rect 797 181 867 197
rect 797 147 813 181
rect 851 147 867 181
rect 797 100 867 147
rect 925 181 995 197
rect 925 147 941 181
rect 979 147 995 181
rect 925 100 995 147
rect 1053 181 1123 197
rect 1053 147 1069 181
rect 1107 147 1123 181
rect 1053 100 1123 147
rect 1181 181 1251 197
rect 1181 147 1197 181
rect 1235 147 1251 181
rect 1181 100 1251 147
rect 1309 181 1379 197
rect 1309 147 1325 181
rect 1363 147 1379 181
rect 1309 100 1379 147
rect 1437 181 1507 197
rect 1437 147 1453 181
rect 1491 147 1507 181
rect 1437 100 1507 147
rect 1565 181 1635 197
rect 1565 147 1581 181
rect 1619 147 1635 181
rect 1565 100 1635 147
rect 1693 181 1763 197
rect 1693 147 1709 181
rect 1747 147 1763 181
rect 1693 100 1763 147
rect 1821 181 1891 197
rect 1821 147 1837 181
rect 1875 147 1891 181
rect 1821 100 1891 147
rect -1891 -147 -1821 -100
rect -1891 -181 -1875 -147
rect -1837 -181 -1821 -147
rect -1891 -197 -1821 -181
rect -1763 -147 -1693 -100
rect -1763 -181 -1747 -147
rect -1709 -181 -1693 -147
rect -1763 -197 -1693 -181
rect -1635 -147 -1565 -100
rect -1635 -181 -1619 -147
rect -1581 -181 -1565 -147
rect -1635 -197 -1565 -181
rect -1507 -147 -1437 -100
rect -1507 -181 -1491 -147
rect -1453 -181 -1437 -147
rect -1507 -197 -1437 -181
rect -1379 -147 -1309 -100
rect -1379 -181 -1363 -147
rect -1325 -181 -1309 -147
rect -1379 -197 -1309 -181
rect -1251 -147 -1181 -100
rect -1251 -181 -1235 -147
rect -1197 -181 -1181 -147
rect -1251 -197 -1181 -181
rect -1123 -147 -1053 -100
rect -1123 -181 -1107 -147
rect -1069 -181 -1053 -147
rect -1123 -197 -1053 -181
rect -995 -147 -925 -100
rect -995 -181 -979 -147
rect -941 -181 -925 -147
rect -995 -197 -925 -181
rect -867 -147 -797 -100
rect -867 -181 -851 -147
rect -813 -181 -797 -147
rect -867 -197 -797 -181
rect -739 -147 -669 -100
rect -739 -181 -723 -147
rect -685 -181 -669 -147
rect -739 -197 -669 -181
rect -611 -147 -541 -100
rect -611 -181 -595 -147
rect -557 -181 -541 -147
rect -611 -197 -541 -181
rect -483 -147 -413 -100
rect -483 -181 -467 -147
rect -429 -181 -413 -147
rect -483 -197 -413 -181
rect -355 -147 -285 -100
rect -355 -181 -339 -147
rect -301 -181 -285 -147
rect -355 -197 -285 -181
rect -227 -147 -157 -100
rect -227 -181 -211 -147
rect -173 -181 -157 -147
rect -227 -197 -157 -181
rect -99 -147 -29 -100
rect -99 -181 -83 -147
rect -45 -181 -29 -147
rect -99 -197 -29 -181
rect 29 -147 99 -100
rect 29 -181 45 -147
rect 83 -181 99 -147
rect 29 -197 99 -181
rect 157 -147 227 -100
rect 157 -181 173 -147
rect 211 -181 227 -147
rect 157 -197 227 -181
rect 285 -147 355 -100
rect 285 -181 301 -147
rect 339 -181 355 -147
rect 285 -197 355 -181
rect 413 -147 483 -100
rect 413 -181 429 -147
rect 467 -181 483 -147
rect 413 -197 483 -181
rect 541 -147 611 -100
rect 541 -181 557 -147
rect 595 -181 611 -147
rect 541 -197 611 -181
rect 669 -147 739 -100
rect 669 -181 685 -147
rect 723 -181 739 -147
rect 669 -197 739 -181
rect 797 -147 867 -100
rect 797 -181 813 -147
rect 851 -181 867 -147
rect 797 -197 867 -181
rect 925 -147 995 -100
rect 925 -181 941 -147
rect 979 -181 995 -147
rect 925 -197 995 -181
rect 1053 -147 1123 -100
rect 1053 -181 1069 -147
rect 1107 -181 1123 -147
rect 1053 -197 1123 -181
rect 1181 -147 1251 -100
rect 1181 -181 1197 -147
rect 1235 -181 1251 -147
rect 1181 -197 1251 -181
rect 1309 -147 1379 -100
rect 1309 -181 1325 -147
rect 1363 -181 1379 -147
rect 1309 -197 1379 -181
rect 1437 -147 1507 -100
rect 1437 -181 1453 -147
rect 1491 -181 1507 -147
rect 1437 -197 1507 -181
rect 1565 -147 1635 -100
rect 1565 -181 1581 -147
rect 1619 -181 1635 -147
rect 1565 -197 1635 -181
rect 1693 -147 1763 -100
rect 1693 -181 1709 -147
rect 1747 -181 1763 -147
rect 1693 -197 1763 -181
rect 1821 -147 1891 -100
rect 1821 -181 1837 -147
rect 1875 -181 1891 -147
rect 1821 -197 1891 -181
<< polycont >>
rect -1875 147 -1837 181
rect -1747 147 -1709 181
rect -1619 147 -1581 181
rect -1491 147 -1453 181
rect -1363 147 -1325 181
rect -1235 147 -1197 181
rect -1107 147 -1069 181
rect -979 147 -941 181
rect -851 147 -813 181
rect -723 147 -685 181
rect -595 147 -557 181
rect -467 147 -429 181
rect -339 147 -301 181
rect -211 147 -173 181
rect -83 147 -45 181
rect 45 147 83 181
rect 173 147 211 181
rect 301 147 339 181
rect 429 147 467 181
rect 557 147 595 181
rect 685 147 723 181
rect 813 147 851 181
rect 941 147 979 181
rect 1069 147 1107 181
rect 1197 147 1235 181
rect 1325 147 1363 181
rect 1453 147 1491 181
rect 1581 147 1619 181
rect 1709 147 1747 181
rect 1837 147 1875 181
rect -1875 -181 -1837 -147
rect -1747 -181 -1709 -147
rect -1619 -181 -1581 -147
rect -1491 -181 -1453 -147
rect -1363 -181 -1325 -147
rect -1235 -181 -1197 -147
rect -1107 -181 -1069 -147
rect -979 -181 -941 -147
rect -851 -181 -813 -147
rect -723 -181 -685 -147
rect -595 -181 -557 -147
rect -467 -181 -429 -147
rect -339 -181 -301 -147
rect -211 -181 -173 -147
rect -83 -181 -45 -147
rect 45 -181 83 -147
rect 173 -181 211 -147
rect 301 -181 339 -147
rect 429 -181 467 -147
rect 557 -181 595 -147
rect 685 -181 723 -147
rect 813 -181 851 -147
rect 941 -181 979 -147
rect 1069 -181 1107 -147
rect 1197 -181 1235 -147
rect 1325 -181 1363 -147
rect 1453 -181 1491 -147
rect 1581 -181 1619 -147
rect 1709 -181 1747 -147
rect 1837 -181 1875 -147
<< locali >>
rect -2051 249 -1955 283
rect 1955 249 2051 283
rect -2051 187 -2017 249
rect 2017 187 2051 249
rect -1891 147 -1875 181
rect -1837 147 -1821 181
rect -1763 147 -1747 181
rect -1709 147 -1693 181
rect -1635 147 -1619 181
rect -1581 147 -1565 181
rect -1507 147 -1491 181
rect -1453 147 -1437 181
rect -1379 147 -1363 181
rect -1325 147 -1309 181
rect -1251 147 -1235 181
rect -1197 147 -1181 181
rect -1123 147 -1107 181
rect -1069 147 -1053 181
rect -995 147 -979 181
rect -941 147 -925 181
rect -867 147 -851 181
rect -813 147 -797 181
rect -739 147 -723 181
rect -685 147 -669 181
rect -611 147 -595 181
rect -557 147 -541 181
rect -483 147 -467 181
rect -429 147 -413 181
rect -355 147 -339 181
rect -301 147 -285 181
rect -227 147 -211 181
rect -173 147 -157 181
rect -99 147 -83 181
rect -45 147 -29 181
rect 29 147 45 181
rect 83 147 99 181
rect 157 147 173 181
rect 211 147 227 181
rect 285 147 301 181
rect 339 147 355 181
rect 413 147 429 181
rect 467 147 483 181
rect 541 147 557 181
rect 595 147 611 181
rect 669 147 685 181
rect 723 147 739 181
rect 797 147 813 181
rect 851 147 867 181
rect 925 147 941 181
rect 979 147 995 181
rect 1053 147 1069 181
rect 1107 147 1123 181
rect 1181 147 1197 181
rect 1235 147 1251 181
rect 1309 147 1325 181
rect 1363 147 1379 181
rect 1437 147 1453 181
rect 1491 147 1507 181
rect 1565 147 1581 181
rect 1619 147 1635 181
rect 1693 147 1709 181
rect 1747 147 1763 181
rect 1821 147 1837 181
rect 1875 147 1891 181
rect -1937 88 -1903 104
rect -1937 -104 -1903 -88
rect -1809 88 -1775 104
rect -1809 -104 -1775 -88
rect -1681 88 -1647 104
rect -1681 -104 -1647 -88
rect -1553 88 -1519 104
rect -1553 -104 -1519 -88
rect -1425 88 -1391 104
rect -1425 -104 -1391 -88
rect -1297 88 -1263 104
rect -1297 -104 -1263 -88
rect -1169 88 -1135 104
rect -1169 -104 -1135 -88
rect -1041 88 -1007 104
rect -1041 -104 -1007 -88
rect -913 88 -879 104
rect -913 -104 -879 -88
rect -785 88 -751 104
rect -785 -104 -751 -88
rect -657 88 -623 104
rect -657 -104 -623 -88
rect -529 88 -495 104
rect -529 -104 -495 -88
rect -401 88 -367 104
rect -401 -104 -367 -88
rect -273 88 -239 104
rect -273 -104 -239 -88
rect -145 88 -111 104
rect -145 -104 -111 -88
rect -17 88 17 104
rect -17 -104 17 -88
rect 111 88 145 104
rect 111 -104 145 -88
rect 239 88 273 104
rect 239 -104 273 -88
rect 367 88 401 104
rect 367 -104 401 -88
rect 495 88 529 104
rect 495 -104 529 -88
rect 623 88 657 104
rect 623 -104 657 -88
rect 751 88 785 104
rect 751 -104 785 -88
rect 879 88 913 104
rect 879 -104 913 -88
rect 1007 88 1041 104
rect 1007 -104 1041 -88
rect 1135 88 1169 104
rect 1135 -104 1169 -88
rect 1263 88 1297 104
rect 1263 -104 1297 -88
rect 1391 88 1425 104
rect 1391 -104 1425 -88
rect 1519 88 1553 104
rect 1519 -104 1553 -88
rect 1647 88 1681 104
rect 1647 -104 1681 -88
rect 1775 88 1809 104
rect 1775 -104 1809 -88
rect 1903 88 1937 104
rect 1903 -104 1937 -88
rect -1891 -181 -1875 -147
rect -1837 -181 -1821 -147
rect -1763 -181 -1747 -147
rect -1709 -181 -1693 -147
rect -1635 -181 -1619 -147
rect -1581 -181 -1565 -147
rect -1507 -181 -1491 -147
rect -1453 -181 -1437 -147
rect -1379 -181 -1363 -147
rect -1325 -181 -1309 -147
rect -1251 -181 -1235 -147
rect -1197 -181 -1181 -147
rect -1123 -181 -1107 -147
rect -1069 -181 -1053 -147
rect -995 -181 -979 -147
rect -941 -181 -925 -147
rect -867 -181 -851 -147
rect -813 -181 -797 -147
rect -739 -181 -723 -147
rect -685 -181 -669 -147
rect -611 -181 -595 -147
rect -557 -181 -541 -147
rect -483 -181 -467 -147
rect -429 -181 -413 -147
rect -355 -181 -339 -147
rect -301 -181 -285 -147
rect -227 -181 -211 -147
rect -173 -181 -157 -147
rect -99 -181 -83 -147
rect -45 -181 -29 -147
rect 29 -181 45 -147
rect 83 -181 99 -147
rect 157 -181 173 -147
rect 211 -181 227 -147
rect 285 -181 301 -147
rect 339 -181 355 -147
rect 413 -181 429 -147
rect 467 -181 483 -147
rect 541 -181 557 -147
rect 595 -181 611 -147
rect 669 -181 685 -147
rect 723 -181 739 -147
rect 797 -181 813 -147
rect 851 -181 867 -147
rect 925 -181 941 -147
rect 979 -181 995 -147
rect 1053 -181 1069 -147
rect 1107 -181 1123 -147
rect 1181 -181 1197 -147
rect 1235 -181 1251 -147
rect 1309 -181 1325 -147
rect 1363 -181 1379 -147
rect 1437 -181 1453 -147
rect 1491 -181 1507 -147
rect 1565 -181 1581 -147
rect 1619 -181 1635 -147
rect 1693 -181 1709 -147
rect 1747 -181 1763 -147
rect 1821 -181 1837 -147
rect 1875 -181 1891 -147
rect -2051 -249 -2017 -187
rect 2017 -249 2051 -187
rect -2051 -283 -1955 -249
rect 1955 -283 2051 -249
<< viali >>
rect -1875 147 -1837 181
rect -1747 147 -1709 181
rect -1619 147 -1581 181
rect -1491 147 -1453 181
rect -1363 147 -1325 181
rect -1235 147 -1197 181
rect -1107 147 -1069 181
rect -979 147 -941 181
rect -851 147 -813 181
rect -723 147 -685 181
rect -595 147 -557 181
rect -467 147 -429 181
rect -339 147 -301 181
rect -211 147 -173 181
rect -83 147 -45 181
rect 45 147 83 181
rect 173 147 211 181
rect 301 147 339 181
rect 429 147 467 181
rect 557 147 595 181
rect 685 147 723 181
rect 813 147 851 181
rect 941 147 979 181
rect 1069 147 1107 181
rect 1197 147 1235 181
rect 1325 147 1363 181
rect 1453 147 1491 181
rect 1581 147 1619 181
rect 1709 147 1747 181
rect 1837 147 1875 181
rect -1937 -88 -1903 88
rect -1809 -88 -1775 88
rect -1681 -88 -1647 88
rect -1553 -88 -1519 88
rect -1425 -88 -1391 88
rect -1297 -88 -1263 88
rect -1169 -88 -1135 88
rect -1041 -88 -1007 88
rect -913 -88 -879 88
rect -785 -88 -751 88
rect -657 -88 -623 88
rect -529 -88 -495 88
rect -401 -88 -367 88
rect -273 -88 -239 88
rect -145 -88 -111 88
rect -17 -88 17 88
rect 111 -88 145 88
rect 239 -88 273 88
rect 367 -88 401 88
rect 495 -88 529 88
rect 623 -88 657 88
rect 751 -88 785 88
rect 879 -88 913 88
rect 1007 -88 1041 88
rect 1135 -88 1169 88
rect 1263 -88 1297 88
rect 1391 -88 1425 88
rect 1519 -88 1553 88
rect 1647 -88 1681 88
rect 1775 -88 1809 88
rect 1903 -88 1937 88
rect -1875 -181 -1837 -147
rect -1747 -181 -1709 -147
rect -1619 -181 -1581 -147
rect -1491 -181 -1453 -147
rect -1363 -181 -1325 -147
rect -1235 -181 -1197 -147
rect -1107 -181 -1069 -147
rect -979 -181 -941 -147
rect -851 -181 -813 -147
rect -723 -181 -685 -147
rect -595 -181 -557 -147
rect -467 -181 -429 -147
rect -339 -181 -301 -147
rect -211 -181 -173 -147
rect -83 -181 -45 -147
rect 45 -181 83 -147
rect 173 -181 211 -147
rect 301 -181 339 -147
rect 429 -181 467 -147
rect 557 -181 595 -147
rect 685 -181 723 -147
rect 813 -181 851 -147
rect 941 -181 979 -147
rect 1069 -181 1107 -147
rect 1197 -181 1235 -147
rect 1325 -181 1363 -147
rect 1453 -181 1491 -147
rect 1581 -181 1619 -147
rect 1709 -181 1747 -147
rect 1837 -181 1875 -147
<< metal1 >>
rect -1887 181 -1825 187
rect -1887 147 -1875 181
rect -1837 147 -1825 181
rect -1887 141 -1825 147
rect -1759 181 -1697 187
rect -1759 147 -1747 181
rect -1709 147 -1697 181
rect -1759 141 -1697 147
rect -1631 181 -1569 187
rect -1631 147 -1619 181
rect -1581 147 -1569 181
rect -1631 141 -1569 147
rect -1503 181 -1441 187
rect -1503 147 -1491 181
rect -1453 147 -1441 181
rect -1503 141 -1441 147
rect -1375 181 -1313 187
rect -1375 147 -1363 181
rect -1325 147 -1313 181
rect -1375 141 -1313 147
rect -1247 181 -1185 187
rect -1247 147 -1235 181
rect -1197 147 -1185 181
rect -1247 141 -1185 147
rect -1119 181 -1057 187
rect -1119 147 -1107 181
rect -1069 147 -1057 181
rect -1119 141 -1057 147
rect -991 181 -929 187
rect -991 147 -979 181
rect -941 147 -929 181
rect -991 141 -929 147
rect -863 181 -801 187
rect -863 147 -851 181
rect -813 147 -801 181
rect -863 141 -801 147
rect -735 181 -673 187
rect -735 147 -723 181
rect -685 147 -673 181
rect -735 141 -673 147
rect -607 181 -545 187
rect -607 147 -595 181
rect -557 147 -545 181
rect -607 141 -545 147
rect -479 181 -417 187
rect -479 147 -467 181
rect -429 147 -417 181
rect -479 141 -417 147
rect -351 181 -289 187
rect -351 147 -339 181
rect -301 147 -289 181
rect -351 141 -289 147
rect -223 181 -161 187
rect -223 147 -211 181
rect -173 147 -161 181
rect -223 141 -161 147
rect -95 181 -33 187
rect -95 147 -83 181
rect -45 147 -33 181
rect -95 141 -33 147
rect 33 181 95 187
rect 33 147 45 181
rect 83 147 95 181
rect 33 141 95 147
rect 161 181 223 187
rect 161 147 173 181
rect 211 147 223 181
rect 161 141 223 147
rect 289 181 351 187
rect 289 147 301 181
rect 339 147 351 181
rect 289 141 351 147
rect 417 181 479 187
rect 417 147 429 181
rect 467 147 479 181
rect 417 141 479 147
rect 545 181 607 187
rect 545 147 557 181
rect 595 147 607 181
rect 545 141 607 147
rect 673 181 735 187
rect 673 147 685 181
rect 723 147 735 181
rect 673 141 735 147
rect 801 181 863 187
rect 801 147 813 181
rect 851 147 863 181
rect 801 141 863 147
rect 929 181 991 187
rect 929 147 941 181
rect 979 147 991 181
rect 929 141 991 147
rect 1057 181 1119 187
rect 1057 147 1069 181
rect 1107 147 1119 181
rect 1057 141 1119 147
rect 1185 181 1247 187
rect 1185 147 1197 181
rect 1235 147 1247 181
rect 1185 141 1247 147
rect 1313 181 1375 187
rect 1313 147 1325 181
rect 1363 147 1375 181
rect 1313 141 1375 147
rect 1441 181 1503 187
rect 1441 147 1453 181
rect 1491 147 1503 181
rect 1441 141 1503 147
rect 1569 181 1631 187
rect 1569 147 1581 181
rect 1619 147 1631 181
rect 1569 141 1631 147
rect 1697 181 1759 187
rect 1697 147 1709 181
rect 1747 147 1759 181
rect 1697 141 1759 147
rect 1825 181 1887 187
rect 1825 147 1837 181
rect 1875 147 1887 181
rect 1825 141 1887 147
rect -1943 88 -1897 100
rect -1943 -88 -1937 88
rect -1903 -88 -1897 88
rect -1943 -100 -1897 -88
rect -1815 88 -1769 100
rect -1815 -88 -1809 88
rect -1775 -88 -1769 88
rect -1815 -100 -1769 -88
rect -1687 88 -1641 100
rect -1687 -88 -1681 88
rect -1647 -88 -1641 88
rect -1687 -100 -1641 -88
rect -1559 88 -1513 100
rect -1559 -88 -1553 88
rect -1519 -88 -1513 88
rect -1559 -100 -1513 -88
rect -1431 88 -1385 100
rect -1431 -88 -1425 88
rect -1391 -88 -1385 88
rect -1431 -100 -1385 -88
rect -1303 88 -1257 100
rect -1303 -88 -1297 88
rect -1263 -88 -1257 88
rect -1303 -100 -1257 -88
rect -1175 88 -1129 100
rect -1175 -88 -1169 88
rect -1135 -88 -1129 88
rect -1175 -100 -1129 -88
rect -1047 88 -1001 100
rect -1047 -88 -1041 88
rect -1007 -88 -1001 88
rect -1047 -100 -1001 -88
rect -919 88 -873 100
rect -919 -88 -913 88
rect -879 -88 -873 88
rect -919 -100 -873 -88
rect -791 88 -745 100
rect -791 -88 -785 88
rect -751 -88 -745 88
rect -791 -100 -745 -88
rect -663 88 -617 100
rect -663 -88 -657 88
rect -623 -88 -617 88
rect -663 -100 -617 -88
rect -535 88 -489 100
rect -535 -88 -529 88
rect -495 -88 -489 88
rect -535 -100 -489 -88
rect -407 88 -361 100
rect -407 -88 -401 88
rect -367 -88 -361 88
rect -407 -100 -361 -88
rect -279 88 -233 100
rect -279 -88 -273 88
rect -239 -88 -233 88
rect -279 -100 -233 -88
rect -151 88 -105 100
rect -151 -88 -145 88
rect -111 -88 -105 88
rect -151 -100 -105 -88
rect -23 88 23 100
rect -23 -88 -17 88
rect 17 -88 23 88
rect -23 -100 23 -88
rect 105 88 151 100
rect 105 -88 111 88
rect 145 -88 151 88
rect 105 -100 151 -88
rect 233 88 279 100
rect 233 -88 239 88
rect 273 -88 279 88
rect 233 -100 279 -88
rect 361 88 407 100
rect 361 -88 367 88
rect 401 -88 407 88
rect 361 -100 407 -88
rect 489 88 535 100
rect 489 -88 495 88
rect 529 -88 535 88
rect 489 -100 535 -88
rect 617 88 663 100
rect 617 -88 623 88
rect 657 -88 663 88
rect 617 -100 663 -88
rect 745 88 791 100
rect 745 -88 751 88
rect 785 -88 791 88
rect 745 -100 791 -88
rect 873 88 919 100
rect 873 -88 879 88
rect 913 -88 919 88
rect 873 -100 919 -88
rect 1001 88 1047 100
rect 1001 -88 1007 88
rect 1041 -88 1047 88
rect 1001 -100 1047 -88
rect 1129 88 1175 100
rect 1129 -88 1135 88
rect 1169 -88 1175 88
rect 1129 -100 1175 -88
rect 1257 88 1303 100
rect 1257 -88 1263 88
rect 1297 -88 1303 88
rect 1257 -100 1303 -88
rect 1385 88 1431 100
rect 1385 -88 1391 88
rect 1425 -88 1431 88
rect 1385 -100 1431 -88
rect 1513 88 1559 100
rect 1513 -88 1519 88
rect 1553 -88 1559 88
rect 1513 -100 1559 -88
rect 1641 88 1687 100
rect 1641 -88 1647 88
rect 1681 -88 1687 88
rect 1641 -100 1687 -88
rect 1769 88 1815 100
rect 1769 -88 1775 88
rect 1809 -88 1815 88
rect 1769 -100 1815 -88
rect 1897 88 1943 100
rect 1897 -88 1903 88
rect 1937 -88 1943 88
rect 1897 -100 1943 -88
rect -1887 -147 -1825 -141
rect -1887 -181 -1875 -147
rect -1837 -181 -1825 -147
rect -1887 -187 -1825 -181
rect -1759 -147 -1697 -141
rect -1759 -181 -1747 -147
rect -1709 -181 -1697 -147
rect -1759 -187 -1697 -181
rect -1631 -147 -1569 -141
rect -1631 -181 -1619 -147
rect -1581 -181 -1569 -147
rect -1631 -187 -1569 -181
rect -1503 -147 -1441 -141
rect -1503 -181 -1491 -147
rect -1453 -181 -1441 -147
rect -1503 -187 -1441 -181
rect -1375 -147 -1313 -141
rect -1375 -181 -1363 -147
rect -1325 -181 -1313 -147
rect -1375 -187 -1313 -181
rect -1247 -147 -1185 -141
rect -1247 -181 -1235 -147
rect -1197 -181 -1185 -147
rect -1247 -187 -1185 -181
rect -1119 -147 -1057 -141
rect -1119 -181 -1107 -147
rect -1069 -181 -1057 -147
rect -1119 -187 -1057 -181
rect -991 -147 -929 -141
rect -991 -181 -979 -147
rect -941 -181 -929 -147
rect -991 -187 -929 -181
rect -863 -147 -801 -141
rect -863 -181 -851 -147
rect -813 -181 -801 -147
rect -863 -187 -801 -181
rect -735 -147 -673 -141
rect -735 -181 -723 -147
rect -685 -181 -673 -147
rect -735 -187 -673 -181
rect -607 -147 -545 -141
rect -607 -181 -595 -147
rect -557 -181 -545 -147
rect -607 -187 -545 -181
rect -479 -147 -417 -141
rect -479 -181 -467 -147
rect -429 -181 -417 -147
rect -479 -187 -417 -181
rect -351 -147 -289 -141
rect -351 -181 -339 -147
rect -301 -181 -289 -147
rect -351 -187 -289 -181
rect -223 -147 -161 -141
rect -223 -181 -211 -147
rect -173 -181 -161 -147
rect -223 -187 -161 -181
rect -95 -147 -33 -141
rect -95 -181 -83 -147
rect -45 -181 -33 -147
rect -95 -187 -33 -181
rect 33 -147 95 -141
rect 33 -181 45 -147
rect 83 -181 95 -147
rect 33 -187 95 -181
rect 161 -147 223 -141
rect 161 -181 173 -147
rect 211 -181 223 -147
rect 161 -187 223 -181
rect 289 -147 351 -141
rect 289 -181 301 -147
rect 339 -181 351 -147
rect 289 -187 351 -181
rect 417 -147 479 -141
rect 417 -181 429 -147
rect 467 -181 479 -147
rect 417 -187 479 -181
rect 545 -147 607 -141
rect 545 -181 557 -147
rect 595 -181 607 -147
rect 545 -187 607 -181
rect 673 -147 735 -141
rect 673 -181 685 -147
rect 723 -181 735 -147
rect 673 -187 735 -181
rect 801 -147 863 -141
rect 801 -181 813 -147
rect 851 -181 863 -147
rect 801 -187 863 -181
rect 929 -147 991 -141
rect 929 -181 941 -147
rect 979 -181 991 -147
rect 929 -187 991 -181
rect 1057 -147 1119 -141
rect 1057 -181 1069 -147
rect 1107 -181 1119 -147
rect 1057 -187 1119 -181
rect 1185 -147 1247 -141
rect 1185 -181 1197 -147
rect 1235 -181 1247 -147
rect 1185 -187 1247 -181
rect 1313 -147 1375 -141
rect 1313 -181 1325 -147
rect 1363 -181 1375 -147
rect 1313 -187 1375 -181
rect 1441 -147 1503 -141
rect 1441 -181 1453 -147
rect 1491 -181 1503 -147
rect 1441 -187 1503 -181
rect 1569 -147 1631 -141
rect 1569 -181 1581 -147
rect 1619 -181 1631 -147
rect 1569 -187 1631 -181
rect 1697 -147 1759 -141
rect 1697 -181 1709 -147
rect 1747 -181 1759 -147
rect 1697 -187 1759 -181
rect 1825 -147 1887 -141
rect 1825 -181 1837 -147
rect 1875 -181 1887 -147
rect 1825 -187 1887 -181
<< properties >>
string FIXED_BBOX -2034 -266 2034 266
string gencell sky130_fd_pr__pfet_01v8_lvt
string library sky130
string parameters w 1.0 l 0.35 m 1 nf 30 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.35 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
