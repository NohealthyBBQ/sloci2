magic
tech sky130A
magscale 1 2
timestamp 1663033959
<< metal1 >>
rect 14920 682870 15420 682910
rect 14920 682040 14960 682870
rect 15390 682040 15420 682870
rect 14920 668280 15420 682040
rect 14920 668180 23410 668280
rect 14920 668100 23840 668180
rect 14920 668060 23410 668100
rect 55960 662600 56100 662620
rect 55960 662500 55980 662600
rect 56080 662500 56100 662600
rect 55960 662480 56100 662500
rect 56200 661680 56340 661700
rect 56200 661580 56220 661680
rect 56320 661580 56340 661680
rect 56200 661560 56340 661580
rect 56480 661080 56620 661100
rect 56480 660980 56500 661080
rect 56600 660980 56620 661080
rect 56480 660960 56620 660980
rect 56720 660560 56860 660580
rect 56720 660460 56740 660560
rect 56840 660460 56860 660560
rect 56720 660440 56860 660460
rect 56980 660200 57120 660220
rect 56980 660100 57000 660200
rect 57100 660100 57120 660200
rect 56980 660080 57120 660100
<< via1 >>
rect 14960 682040 15390 682870
rect 55980 662500 56080 662600
rect 56220 661580 56320 661680
rect 56500 660980 56600 661080
rect 56740 660460 56840 660560
rect 57000 660100 57100 660200
<< metal2 >>
rect 14920 682870 15420 682910
rect 14920 682040 14960 682870
rect 15390 682040 15420 682870
rect 14920 681990 15420 682040
rect 23190 671610 25400 671620
rect 23190 671440 23210 671610
rect 23370 671440 25400 671610
rect 23190 671420 25400 671440
rect 55960 662600 56100 662620
rect 55960 662500 55980 662600
rect 56080 662500 56100 662600
rect 55960 335220 56100 662500
rect 56200 661680 56340 661700
rect 56200 661580 56220 661680
rect 56320 661580 56340 661680
rect 56200 378460 56340 661580
rect 56480 661080 56620 661100
rect 56480 660980 56500 661080
rect 56600 660980 56620 661080
rect 56480 421660 56620 660980
rect 56720 660560 56860 660580
rect 56720 660460 56740 660560
rect 56840 660460 56860 660560
rect 56720 466080 56860 660460
rect 56980 660200 57120 660220
rect 56980 660100 57000 660200
rect 57100 660100 57120 660200
rect 56980 508120 57120 660100
rect 238000 591000 246800 592200
rect 238000 582000 239000 591000
rect 246000 582000 246800 591000
rect 238000 580200 246800 582000
rect 246300 579400 246700 580200
rect 56980 507980 57000 508120
rect 57100 507980 57120 508120
rect 56980 507960 57120 507980
rect 56720 465940 56740 466080
rect 56840 465940 56860 466080
rect 56720 465920 56860 465940
rect 56480 421520 56500 421660
rect 56600 421520 56620 421660
rect 56480 421500 56620 421520
rect 56200 378320 56220 378460
rect 56320 378320 56340 378460
rect 56200 378300 56340 378320
rect 55960 335080 55980 335220
rect 56080 335080 56100 335220
rect 55960 335060 56100 335080
<< via2 >>
rect 14960 682040 15390 682870
rect 23210 671440 23370 671610
rect 239000 582000 246000 591000
rect 57000 507980 57100 508120
rect 56740 465940 56840 466080
rect 56500 421520 56600 421660
rect 56220 378320 56320 378460
rect 55980 335080 56080 335220
<< metal3 >>
rect 16194 702300 21194 704800
rect 68194 702300 73194 704800
rect 120194 703200 125194 704800
rect 17070 689360 19380 702300
rect 68470 689480 70760 702300
rect 42500 689440 70760 689480
rect 17070 689330 26050 689360
rect 17070 688210 41870 689330
rect 42500 688410 42560 689440
rect 43180 688410 70760 689440
rect 42500 688360 70760 688410
rect 120000 701000 125200 703200
rect 165594 702300 170594 704800
rect 175894 702300 180894 704800
rect 17070 688200 26050 688210
rect -800 682910 1700 685242
rect -800 682870 15420 682910
rect -800 682040 14960 682870
rect 15390 682040 15420 682870
rect -800 681990 15420 682040
rect -800 680242 1700 681990
rect 40710 680350 41870 688210
rect 40720 679110 41870 680350
rect 40720 677240 41720 677320
rect 40720 676130 40770 677240
rect 41640 676130 41720 677240
rect 40720 676080 41720 676130
rect 23190 671610 23390 671620
rect 23190 671440 23210 671610
rect 23370 671440 23390 671610
rect 23190 669080 23390 671440
rect 23190 668680 23210 669080
rect 23370 668680 23390 669080
rect 23190 668640 23390 668680
rect 310 648642 1780 648730
rect -800 648600 1780 648642
rect -800 647000 80246 648600
rect -800 643842 73000 647000
rect 246 638642 73000 643842
rect -800 635000 73000 638642
rect 79000 635000 80246 647000
rect -800 633842 80246 635000
rect 246 633838 80246 633842
rect 120000 606000 124000 701000
rect 21990 604000 22000 606000
rect 24000 604000 24010 606000
rect 22000 596000 24000 604000
rect 120000 602000 288000 606000
rect 22000 594000 285400 596000
rect 238990 591000 246010 591005
rect 164000 590000 239000 591000
rect 164000 583000 165000 590000
rect 182000 583000 239000 590000
rect 164000 582000 239000 583000
rect 246000 582000 246010 591000
rect 154000 581400 158000 582000
rect 238990 581995 246010 582000
rect 154000 580000 245900 581400
rect 283800 580600 285400 594000
rect 286000 580600 287600 602000
rect -800 564220 1660 564242
rect -800 564080 4430 564220
rect -800 559570 860 564080
rect 4260 559570 4430 564080
rect -800 559442 4430 559570
rect 680 555000 4430 559442
rect 680 554242 1000 555000
rect -800 550000 1000 554242
rect 4000 550000 4430 555000
rect -800 549442 4430 550000
rect 680 549410 4430 549442
rect 260 508120 57120 508140
rect 260 508096 57000 508120
rect -800 507984 57000 508096
rect 260 507980 57000 507984
rect 57100 507980 57120 508120
rect 260 507960 57120 507980
rect 280 466080 56860 466100
rect 280 466056 56740 466080
rect -800 465944 56740 466056
rect 280 465940 56740 465944
rect 56840 465940 56860 466080
rect 280 465920 56860 465940
rect 360 421660 56620 421680
rect 360 421652 56500 421660
rect -800 421540 56500 421652
rect 360 421520 56500 421540
rect 56600 421520 56620 421660
rect 360 421500 56620 421520
rect 400 378460 56340 378480
rect 400 378430 56220 378460
rect -800 378320 56220 378430
rect 56320 378320 56340 378460
rect -800 378318 56340 378320
rect 400 378300 56340 378318
rect 260 335220 56100 335240
rect 260 335208 55980 335220
rect -800 335096 55980 335208
rect 260 335080 55980 335096
rect 56080 335080 56100 335220
rect 260 335060 56100 335080
rect 200 295532 800 295600
rect -800 295420 800 295532
rect 200 295400 800 295420
rect 154000 295400 158000 580000
rect 200 294600 158000 295400
rect 154000 294000 158000 294600
rect 1650 177690 20600 178000
rect 982 177688 20600 177690
rect -800 177600 20600 177688
rect -800 172888 11600 177600
rect 982 172300 11600 172888
rect 20200 172300 20600 177600
rect 982 171900 20600 172300
rect 982 167688 5298 171900
rect -800 162890 5298 167688
rect -800 162888 1660 162890
<< via3 >>
rect 42560 688410 43180 689440
rect 40770 676130 41640 677240
rect 23210 668680 23370 669080
rect 73000 635000 79000 647000
rect 22000 604000 24000 606000
rect 165000 583000 182000 590000
rect 860 559570 4260 564080
rect 1000 550000 4000 555000
rect 11600 172300 20200 177600
<< metal4 >>
rect 165594 703000 170594 704800
rect 175894 703000 180894 704800
rect 42500 689440 43450 689470
rect 42500 688410 42560 689440
rect 43180 688410 43450 689440
rect 42500 677320 43450 688410
rect 40720 677240 43450 677320
rect 40720 676130 40770 677240
rect 41640 676130 43450 677240
rect 40720 676090 43450 676130
rect 40720 676080 43220 676090
rect 60220 676010 65450 676030
rect 56870 675970 65450 676010
rect 56870 675440 60910 675970
rect 65380 675440 65450 675970
rect 56870 675370 65450 675440
rect 23190 669080 23390 669110
rect 23190 668680 23210 669080
rect 23370 668680 23390 669080
rect 23190 608120 23390 668680
rect 26600 633690 28120 662640
rect 72999 647000 79001 647001
rect 72999 635000 73000 647000
rect 79000 635000 79001 647000
rect 72999 634999 79001 635000
rect 26090 633500 28790 633690
rect 26090 631620 26270 633500
rect 28580 631620 28790 633500
rect 26090 631490 28790 631620
rect 32100 620300 39650 620900
rect 32100 614050 32850 620300
rect 38700 614050 39650 620300
rect 32100 613600 39650 614050
rect 21660 606000 25780 608120
rect 21660 604000 22000 606000
rect 24000 604000 25780 606000
rect 21660 603350 25780 604000
rect 690 564080 4450 564270
rect 690 559570 860 564080
rect 4260 559570 4450 564080
rect 690 559400 4450 559570
rect 999 555000 4001 555001
rect 999 550000 1000 555000
rect 4000 550000 4001 555000
rect 999 549999 4001 550000
rect 30150 178000 39650 613600
rect 165000 590001 182000 703000
rect 305500 645000 316500 646500
rect 164999 590000 182001 590001
rect 164999 583000 165000 590000
rect 182000 583000 182001 590000
rect 164999 582999 182001 583000
rect 238000 584000 248000 636000
rect 305500 637000 307000 645000
rect 315000 637000 316500 645000
rect 238000 580000 260000 584000
rect 305500 580300 316500 637000
rect 238200 570900 240100 574000
rect 258800 571400 260000 580000
rect 238200 568100 239300 570900
rect 238200 563700 240200 568100
rect 239700 558000 240200 563700
rect 510000 563000 526000 660000
rect 263600 557900 316600 558100
rect 510000 555000 511000 563000
rect 525000 555000 526000 563000
rect 510000 554000 526000 555000
rect 11100 177600 39650 178000
rect 11100 172300 11600 177600
rect 20200 172300 39650 177600
rect 11100 171950 39650 172300
rect 11100 171900 34150 171950
<< via4 >>
rect 60910 675440 65380 675970
rect 73000 635000 79000 647000
rect 26270 631620 28580 633500
rect 32850 614050 38700 620300
rect 860 559570 4260 564080
rect 1000 550000 4000 555000
rect 238000 636000 248000 644000
rect 307000 637000 315000 645000
rect 238200 558000 239700 563700
rect 263600 556400 316600 557900
rect 511000 555000 525000 563000
<< metal5 >>
rect 165594 702300 170594 704800
rect 175894 702300 180894 704800
rect 60790 675970 65590 676060
rect 60790 675440 60910 675970
rect 65380 675440 65590 675970
rect 26080 633500 28810 633710
rect 26080 631620 26270 633500
rect 28580 631620 28810 633500
rect 26080 564330 28810 631620
rect 33890 625850 34330 675040
rect 39240 625850 39680 674940
rect 42370 625850 42840 674830
rect 44740 625850 45180 675000
rect 45790 625850 46240 663160
rect 60790 652300 65590 675440
rect 32150 620300 51000 625850
rect 32150 614050 32850 620300
rect 38700 614050 51000 620300
rect 32150 613550 51000 614050
rect 60820 564330 65590 652300
rect 72976 647000 79024 647024
rect 72976 635000 73000 647000
rect 79000 645000 553600 647000
rect 79000 644000 307000 645000
rect 79000 636000 238000 644000
rect 248000 637000 307000 644000
rect 315000 637000 553600 645000
rect 248000 636000 553600 637000
rect 79000 635000 553600 636000
rect 72976 634976 79024 635000
rect 26080 564320 65590 564330
rect 1770 564270 65590 564320
rect 690 564080 65590 564270
rect 690 559570 860 564080
rect 4260 564000 65590 564080
rect 4260 563700 526000 564000
rect 4260 559570 238200 563700
rect 690 559400 238200 559570
rect 1000 558000 238200 559400
rect 239700 563000 526000 563700
rect 239700 558000 511000 563000
rect 1000 557900 511000 558000
rect 1000 556400 263600 557900
rect 316600 556400 511000 557900
rect 1000 555024 511000 556400
rect 976 555000 511000 555024
rect 525000 555000 526000 563000
rect 976 550000 1000 555000
rect 4000 550000 526000 555000
rect 976 549976 4024 550000
<< comment >>
rect -100 704000 584100 704100
rect -100 0 0 704000
rect 584000 0 584100 704000
rect -100 -100 584100 0
use BGR_lvs  BGR_lvs_0
timestamp 1663029885
transform 1 0 254230 0 1 568403
box -14230 -10403 62405 12600
use VCO  VCO_0
timestamp 1663030914
transform 1 0 -7837 0 1 638742
box 31141 20430 65400 41673
<< labels >>
flabel metal3 s -800 295420 480 295532 0 FreeSans 1120 0 0 0 gpio_analog[12]
port 3 nsew signal bidirectional
flabel metal3 0 680242 1700 685242 0 FreeSans 1120 0 0 0 io_analog[10]
flabel metal3 s 175894 702300 180894 704800 0 FreeSans 1920 180 0 0 io_analog[6]
port 43 nsew signal bidirectional
flabel metal4 s 175894 702300 180894 704800 0 FreeSans 1920 180 0 0 io_analog[6]
port 43 nsew signal bidirectional
flabel metal5 s 175894 702300 180894 704800 0 FreeSans 1920 180 0 0 io_analog[6]
port 43 nsew signal bidirectional
flabel metal3 s 120194 702300 125194 704800 0 FreeSans 1920 180 0 0 io_analog[7]
port 44 nsew signal bidirectional
flabel metal3 s 68194 702300 73194 704800 0 FreeSans 1920 180 0 0 io_analog[8]
port 45 nsew signal bidirectional
flabel metal3 s 16194 702300 21194 704800 0 FreeSans 1920 180 0 0 io_analog[9]
port 46 nsew signal bidirectional
flabel metal3 s 165594 702300 170594 704800 0 FreeSans 1920 180 0 0 io_analog[6]
port 49 nsew signal bidirectional
flabel metal4 s 165594 702300 170594 704800 0 FreeSans 1920 180 0 0 io_analog[6]
port 49 nsew signal bidirectional
flabel metal5 s 165594 702300 170594 704800 0 FreeSans 1920 180 0 0 io_analog[6]
port 49 nsew signal bidirectional
flabel metal3 s -800 507984 480 508096 0 FreeSans 1120 0 0 0 io_in[14]
port 61 nsew signal input
flabel metal3 s -800 421540 480 421652 0 FreeSans 1120 0 0 0 io_in[16]
port 63 nsew signal input
flabel metal3 s -800 378318 480 378430 0 FreeSans 1120 0 0 0 io_in[17]
port 64 nsew signal input
flabel metal3 s -800 335096 480 335208 0 FreeSans 1120 0 0 0 io_in[18]
port 65 nsew signal input
flabel metal3 s -800 465944 480 466056 0 FreeSans 1120 0 0 0 io_in_3v3[15]
port 89 nsew signal input
flabel metal3 s 0 643842 1660 648642 0 FreeSans 1120 0 0 0 vccd2
port 554 nsew signal bidirectional
flabel metal3 s 0 633842 1660 638642 0 FreeSans 1120 0 0 0 vccd2
port 555 nsew signal bidirectional
flabel metal3 s 0 559442 1660 564242 0 FreeSans 1120 0 0 0 vssa2
port 566 nsew signal bidirectional
flabel metal3 s 0 549442 1660 554242 0 FreeSans 1120 0 0 0 vssa2
port 567 nsew signal bidirectional
flabel metal3 s 0 172888 1660 177688 0 FreeSans 1120 0 0 0 vssd2
port 570 nsew signal bidirectional
flabel metal3 s 0 162888 1660 167688 0 FreeSans 1120 0 0 0 vssd2
port 571 nsew signal bidirectional
flabel metal5 26080 559400 65590 564330 0 FreeSans 16000 0 0 0 GND
rlabel metal2 56980 508120 57120 660100 1 CTRL1
rlabel metal2 56720 466080 56860 660460 1 CTRL2
rlabel metal2 56480 421660 56620 660980 1 CTRL3
rlabel metal2 56200 378460 56340 661580 1 CTRL4
rlabel metal2 55960 335220 56100 662500 1 CTRL5
flabel metal1 14920 668060 15420 682040 0 FreeSans 8000 0 0 0 VCTRL
flabel metal4 21660 603350 25780 608120 0 FreeSans 8000 0 0 0 REF
rlabel metal3 17070 688210 41870 689330 1 OUT0
rlabel metal3 43180 688360 70760 689480 1 OUT180
<< properties >>
string FIXED_BBOX 0 0 584000 704000
<< end >>
