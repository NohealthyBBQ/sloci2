magic
tech sky130A
magscale 1 2
timestamp 1662665484
<< nwell >>
rect 17100 7240 19040 7245
rect 17710 5070 19040 7240
rect 17710 4990 17780 5070
rect 18360 4990 18420 5070
rect 18620 5020 19040 5070
rect 19035 4990 19040 5020
rect 18180 4384 18600 4390
rect 17930 210 18350 4384
rect 20550 2400 20750 5650
<< locali >>
rect 17670 7175 17825 7215
rect 18315 7170 18470 7210
rect 18970 6975 20025 7020
rect 19990 6180 20025 6975
rect 20520 5545 20775 5580
rect 17535 4310 17570 5060
rect 17670 5030 17825 5070
rect 18070 4350 18105 5060
rect 18185 4350 18220 5060
rect 18320 5030 18475 5070
rect 18070 4315 18220 4350
rect 18715 4315 18750 5065
rect 18185 4310 18220 4315
rect 19075 4105 19110 4270
rect 19870 4105 19905 4270
rect 20735 4070 20770 4075
rect 19985 3930 20020 4070
rect 20515 4035 20775 4070
rect 20520 3980 20555 4035
rect 20735 3980 20770 4035
rect 20510 3935 20770 3980
rect 21265 3940 21300 4080
rect 20515 2435 20770 2470
rect 18070 245 18220 280
rect 18070 -100 18220 -65
rect 19070 -100 19115 790
rect 19370 -95 19410 780
rect 18070 -615 18220 -580
<< metal1 >>
rect 17220 7150 20470 7220
rect 17220 5180 17280 7150
rect 17310 7110 17400 7120
rect 17310 7050 17320 7110
rect 17390 7100 17400 7110
rect 17390 7050 17530 7100
rect 17310 7040 17400 7050
rect 17440 6980 17530 6990
rect 17440 6970 17450 6980
rect 17310 6920 17450 6970
rect 17520 6920 17530 6980
rect 17440 6910 17530 6920
rect 17310 6850 17400 6860
rect 17310 6790 17320 6850
rect 17390 6840 17400 6850
rect 17390 6790 17530 6840
rect 17310 6780 17400 6790
rect 17440 6720 17530 6730
rect 17310 6670 17450 6720
rect 17440 6660 17450 6670
rect 17520 6660 17530 6720
rect 17440 6650 17530 6660
rect 17310 6590 17400 6600
rect 17310 6530 17320 6590
rect 17390 6540 17530 6590
rect 17390 6530 17400 6540
rect 17310 6520 17400 6530
rect 17440 6460 17530 6470
rect 17310 6410 17450 6460
rect 17440 6400 17450 6410
rect 17520 6400 17530 6460
rect 17440 6390 17530 6400
rect 17310 6330 17400 6340
rect 17310 6270 17320 6330
rect 17390 6280 17530 6330
rect 17390 6270 17400 6280
rect 17310 6260 17400 6270
rect 17440 6210 17530 6220
rect 17440 6200 17450 6210
rect 17310 6160 17450 6200
rect 17440 6150 17450 6160
rect 17520 6150 17530 6210
rect 17440 6140 17530 6150
rect 17310 6080 17400 6090
rect 17310 6020 17320 6080
rect 17390 6030 17530 6080
rect 17390 6020 17400 6030
rect 17310 6010 17400 6020
rect 17440 5960 17530 5970
rect 17440 5950 17450 5960
rect 17310 5900 17450 5950
rect 17520 5900 17530 5960
rect 17440 5890 17530 5900
rect 17310 5830 17400 5840
rect 17310 5770 17320 5830
rect 17390 5820 17400 5830
rect 17390 5770 17530 5820
rect 17310 5760 17400 5770
rect 17440 5700 17530 5710
rect 17440 5690 17450 5700
rect 17310 5640 17450 5690
rect 17520 5640 17530 5700
rect 17440 5630 17530 5640
rect 17310 5570 17400 5580
rect 17310 5510 17320 5570
rect 17390 5560 17400 5570
rect 17390 5520 17530 5560
rect 17390 5510 17400 5520
rect 17310 5500 17400 5510
rect 17440 5440 17530 5450
rect 17310 5390 17450 5440
rect 17440 5380 17450 5390
rect 17520 5380 17530 5440
rect 17440 5370 17530 5380
rect 17310 5310 17400 5320
rect 17310 5250 17320 5310
rect 17390 5260 17530 5310
rect 17390 5250 17400 5260
rect 17310 5240 17400 5250
rect 17440 5180 17530 5190
rect 17560 5180 17620 7150
rect 17870 5180 17930 7150
rect 17960 7110 18050 7120
rect 17960 7050 17970 7110
rect 18040 7100 18050 7110
rect 18040 7050 18180 7100
rect 17960 7040 18050 7050
rect 18090 6980 18180 6990
rect 18090 6972 18100 6980
rect 17969 6970 18100 6972
rect 17960 6920 18100 6970
rect 18170 6920 18180 6980
rect 18090 6910 18180 6920
rect 17960 6850 18050 6860
rect 17960 6790 17970 6850
rect 18040 6844 18050 6850
rect 18040 6840 18169 6844
rect 18040 6790 18180 6840
rect 17960 6780 18050 6790
rect 18090 6720 18180 6730
rect 17960 6670 18100 6720
rect 18090 6660 18100 6670
rect 18170 6660 18180 6720
rect 18090 6650 18180 6660
rect 17960 6590 18050 6600
rect 17960 6530 17970 6590
rect 18040 6540 18180 6590
rect 18040 6530 18050 6540
rect 17960 6520 18050 6530
rect 18090 6460 18180 6470
rect 17960 6410 18100 6460
rect 18090 6400 18100 6410
rect 18170 6400 18180 6460
rect 18090 6390 18180 6400
rect 17960 6332 18050 6340
rect 17960 6330 18169 6332
rect 17960 6270 17970 6330
rect 18040 6280 18180 6330
rect 18040 6270 18050 6280
rect 17960 6260 18050 6270
rect 18090 6210 18180 6220
rect 18090 6204 18100 6210
rect 17969 6200 18100 6204
rect 17960 6160 18100 6200
rect 17969 6158 18100 6160
rect 18090 6150 18100 6158
rect 18170 6150 18180 6210
rect 18090 6140 18180 6150
rect 17960 6080 18050 6090
rect 17960 6020 17970 6080
rect 18040 6030 18180 6080
rect 18040 6020 18050 6030
rect 17960 6010 18050 6020
rect 18090 5960 18180 5970
rect 18090 5950 18100 5960
rect 17960 5900 18100 5950
rect 18170 5900 18180 5960
rect 18090 5890 18180 5900
rect 17960 5830 18050 5840
rect 17960 5770 17970 5830
rect 18040 5820 18050 5830
rect 18040 5770 18180 5820
rect 17960 5760 18050 5770
rect 18090 5700 18180 5710
rect 18090 5692 18100 5700
rect 17969 5690 18100 5692
rect 17960 5640 18100 5690
rect 18170 5640 18180 5700
rect 18090 5630 18180 5640
rect 17960 5570 18050 5580
rect 17960 5510 17970 5570
rect 18040 5564 18050 5570
rect 18040 5560 18169 5564
rect 18040 5520 18180 5560
rect 18040 5518 18169 5520
rect 18040 5510 18050 5518
rect 17960 5500 18050 5510
rect 18090 5440 18180 5450
rect 17960 5390 18100 5440
rect 18090 5380 18100 5390
rect 18170 5380 18180 5440
rect 18090 5370 18180 5380
rect 17960 5310 18050 5320
rect 17960 5250 17970 5310
rect 18040 5260 18180 5310
rect 18040 5250 18050 5260
rect 17960 5240 18050 5250
rect 18090 5180 18180 5190
rect 18210 5180 18270 7150
rect 18520 5180 18580 7150
rect 18610 7110 18700 7120
rect 18610 7050 18620 7110
rect 18690 7100 18700 7110
rect 18690 7050 18830 7100
rect 18610 7040 18700 7050
rect 18740 6980 18830 6990
rect 18740 6972 18750 6980
rect 18619 6970 18750 6972
rect 18610 6920 18750 6970
rect 18820 6920 18830 6980
rect 18740 6910 18830 6920
rect 18610 6850 18700 6860
rect 18610 6790 18620 6850
rect 18690 6844 18700 6850
rect 18690 6840 18819 6844
rect 18690 6790 18830 6840
rect 18610 6780 18700 6790
rect 18740 6720 18830 6730
rect 18610 6670 18750 6720
rect 18740 6660 18750 6670
rect 18820 6660 18830 6720
rect 18740 6650 18830 6660
rect 18610 6590 18700 6600
rect 18610 6530 18620 6590
rect 18690 6540 18830 6590
rect 18690 6530 18700 6540
rect 18610 6520 18700 6530
rect 18740 6460 18830 6470
rect 18610 6410 18750 6460
rect 18740 6400 18750 6410
rect 18820 6400 18830 6460
rect 18740 6390 18830 6400
rect 18610 6332 18700 6340
rect 18610 6330 18819 6332
rect 18610 6270 18620 6330
rect 18690 6280 18830 6330
rect 18690 6270 18700 6280
rect 18610 6260 18700 6270
rect 18740 6210 18830 6220
rect 18740 6204 18750 6210
rect 18619 6200 18750 6204
rect 18610 6160 18750 6200
rect 18619 6158 18750 6160
rect 18740 6150 18750 6158
rect 18820 6150 18830 6210
rect 18740 6140 18830 6150
rect 18610 6080 18700 6090
rect 18610 6020 18620 6080
rect 18690 6030 18830 6080
rect 18690 6020 18700 6030
rect 18610 6010 18700 6020
rect 18740 5960 18830 5970
rect 18740 5950 18750 5960
rect 18610 5900 18750 5950
rect 18820 5900 18830 5960
rect 18740 5890 18830 5900
rect 18610 5830 18700 5840
rect 18610 5770 18620 5830
rect 18690 5820 18700 5830
rect 18690 5770 18830 5820
rect 18610 5760 18700 5770
rect 18740 5700 18830 5710
rect 18740 5692 18750 5700
rect 18619 5690 18750 5692
rect 18610 5640 18750 5690
rect 18820 5640 18830 5700
rect 18740 5630 18830 5640
rect 18610 5570 18700 5580
rect 18610 5510 18620 5570
rect 18690 5564 18700 5570
rect 18690 5560 18819 5564
rect 18690 5520 18830 5560
rect 18690 5518 18819 5520
rect 18690 5510 18700 5518
rect 18610 5500 18700 5510
rect 18740 5440 18830 5450
rect 18610 5390 18750 5440
rect 18740 5380 18750 5390
rect 18820 5380 18830 5440
rect 18740 5370 18830 5380
rect 18610 5310 18700 5320
rect 18610 5250 18620 5310
rect 18690 5260 18830 5310
rect 18690 5250 18700 5260
rect 18610 5240 18700 5250
rect 18740 5180 18830 5190
rect 18860 5180 18920 7150
rect 20410 6220 20470 7150
rect 20070 6160 20470 6220
rect 17310 5130 17450 5180
rect 17440 5120 17450 5130
rect 17520 5120 17530 5180
rect 17960 5130 18100 5180
rect 17440 5110 17530 5120
rect 18090 5120 18100 5130
rect 18170 5120 18180 5180
rect 18610 5130 18750 5180
rect 18090 5110 18180 5120
rect 18740 5120 18750 5130
rect 18820 5120 18830 5180
rect 18740 5110 18830 5120
rect 17100 4310 18020 4370
rect 17620 400 17680 4310
rect 17710 4250 17790 4260
rect 17710 4180 17720 4250
rect 17780 4180 17790 4250
rect 17860 4190 17930 4240
rect 17710 4170 17790 4180
rect 17850 4120 17930 4130
rect 17850 4110 17860 4120
rect 17710 4060 17860 4110
rect 17850 4050 17860 4060
rect 17920 4050 17930 4120
rect 17850 4040 17930 4050
rect 17710 3990 17790 4000
rect 17710 3920 17720 3990
rect 17780 3940 17930 3990
rect 17780 3920 17790 3940
rect 17710 3910 17790 3920
rect 17850 3870 17930 3880
rect 17850 3860 17860 3870
rect 17710 3810 17860 3860
rect 17850 3800 17860 3810
rect 17920 3800 17930 3870
rect 17850 3790 17930 3800
rect 17710 3740 17790 3750
rect 17710 3670 17720 3740
rect 17780 3730 17790 3740
rect 17780 3680 17930 3730
rect 17780 3670 17790 3680
rect 17710 3660 17790 3670
rect 17850 3610 17930 3620
rect 17850 3600 17860 3610
rect 17710 3550 17860 3600
rect 17850 3540 17860 3550
rect 17920 3540 17930 3610
rect 17850 3530 17930 3540
rect 17710 3480 17790 3490
rect 17710 3410 17720 3480
rect 17780 3470 17790 3480
rect 17780 3420 17930 3470
rect 17780 3410 17790 3420
rect 17710 3400 17790 3410
rect 17850 3360 17930 3370
rect 17850 3350 17860 3360
rect 17710 3300 17860 3350
rect 17850 3290 17860 3300
rect 17920 3290 17930 3360
rect 17850 3280 17930 3290
rect 17710 3230 17790 3240
rect 17710 3160 17720 3230
rect 17780 3220 17790 3230
rect 17780 3170 17930 3220
rect 17780 3160 17790 3170
rect 17710 3150 17790 3160
rect 17850 3100 17930 3110
rect 17850 3090 17860 3100
rect 17710 3040 17860 3090
rect 17850 3030 17860 3040
rect 17920 3030 17930 3100
rect 17850 3020 17930 3030
rect 17710 2970 17790 2980
rect 17710 2900 17720 2970
rect 17780 2960 17790 2970
rect 17780 2910 17930 2960
rect 17780 2900 17790 2910
rect 17710 2890 17790 2900
rect 17850 2840 17930 2850
rect 17850 2830 17860 2840
rect 17710 2780 17860 2830
rect 17850 2770 17860 2780
rect 17920 2770 17930 2840
rect 17850 2760 17930 2770
rect 17710 2720 17790 2730
rect 17710 2650 17720 2720
rect 17780 2710 17790 2720
rect 17780 2650 17930 2710
rect 17710 2640 17790 2650
rect 17850 2590 17930 2600
rect 17850 2580 17860 2590
rect 17710 2530 17860 2580
rect 17850 2520 17860 2530
rect 17920 2520 17930 2590
rect 17850 2510 17930 2520
rect 17710 2460 17790 2470
rect 17710 2390 17720 2460
rect 17780 2450 17790 2460
rect 17780 2400 17930 2450
rect 17780 2390 17790 2400
rect 17710 2380 17790 2390
rect 17850 2330 17930 2340
rect 17850 2320 17860 2330
rect 17710 2270 17860 2320
rect 17850 2260 17860 2270
rect 17920 2260 17930 2330
rect 17850 2250 17930 2260
rect 17710 2200 17790 2210
rect 17710 2130 17720 2200
rect 17780 2140 17930 2200
rect 17780 2130 17790 2140
rect 17710 2120 17790 2130
rect 17850 2080 17930 2090
rect 17850 2070 17860 2080
rect 17710 2010 17860 2070
rect 17920 2010 17930 2080
rect 17850 2000 17930 2010
rect 17710 1950 17790 1960
rect 17710 1880 17720 1950
rect 17780 1940 17790 1950
rect 17780 1890 17930 1940
rect 17780 1880 17790 1890
rect 17710 1870 17790 1880
rect 17850 1820 17930 1830
rect 17850 1810 17860 1820
rect 17710 1760 17860 1810
rect 17850 1750 17860 1760
rect 17920 1750 17930 1820
rect 17850 1740 17930 1750
rect 17710 1690 17790 1700
rect 17710 1620 17720 1690
rect 17780 1680 17790 1690
rect 17780 1630 17930 1680
rect 17780 1620 17790 1630
rect 17710 1610 17790 1620
rect 17850 1560 17930 1570
rect 17850 1550 17860 1560
rect 17710 1510 17860 1550
rect 17850 1490 17860 1510
rect 17920 1490 17930 1560
rect 17850 1480 17930 1490
rect 17710 1430 17790 1440
rect 17710 1360 17720 1430
rect 17780 1380 17930 1430
rect 17780 1360 17790 1380
rect 17710 1350 17790 1360
rect 17850 1310 17930 1320
rect 17850 1300 17860 1310
rect 17710 1250 17860 1300
rect 17850 1240 17860 1250
rect 17920 1240 17930 1310
rect 17850 1230 17930 1240
rect 17710 1180 17790 1190
rect 17710 1110 17720 1180
rect 17780 1170 17790 1180
rect 17780 1120 17930 1170
rect 17780 1110 17790 1120
rect 17710 1100 17790 1110
rect 17850 1050 17930 1060
rect 17850 1040 17860 1050
rect 17710 990 17860 1040
rect 17850 980 17860 990
rect 17920 980 17930 1050
rect 17850 970 17930 980
rect 17710 920 17790 930
rect 17710 850 17720 920
rect 17780 910 17790 920
rect 17780 860 17930 910
rect 17780 850 17790 860
rect 17710 840 17790 850
rect 17850 800 17930 810
rect 17850 790 17860 800
rect 17710 730 17860 790
rect 17920 730 17930 800
rect 17850 720 17930 730
rect 17710 670 17790 680
rect 17710 600 17720 670
rect 17780 660 17790 670
rect 17780 610 17930 660
rect 17780 600 17790 610
rect 17710 590 17790 600
rect 17850 540 17930 550
rect 17850 530 17860 540
rect 17710 480 17860 530
rect 17850 470 17860 480
rect 17920 470 17930 540
rect 17850 460 17930 470
rect 17710 410 17790 420
rect 17710 340 17720 410
rect 17780 400 17790 410
rect 17960 400 18020 4310
rect 18270 4310 18670 4370
rect 18270 400 18330 4310
rect 18500 4250 18580 4260
rect 18500 4240 18510 4250
rect 18360 4234 18510 4240
rect 18360 4200 18430 4234
rect 18500 4200 18510 4234
rect 18360 4194 18510 4200
rect 18360 4190 18430 4194
rect 18500 4180 18510 4194
rect 18570 4180 18580 4250
rect 18500 4170 18580 4180
rect 18360 4120 18440 4130
rect 18360 4050 18370 4120
rect 18430 4112 18440 4120
rect 18430 4110 18571 4112
rect 18430 4060 18580 4110
rect 18430 4050 18440 4060
rect 18360 4040 18440 4050
rect 18500 3990 18580 4000
rect 18360 3940 18510 3990
rect 18371 3938 18510 3940
rect 18500 3920 18510 3938
rect 18570 3920 18580 3990
rect 18500 3910 18580 3920
rect 18360 3870 18440 3880
rect 18360 3800 18370 3870
rect 18430 3860 18440 3870
rect 18430 3810 18580 3860
rect 18430 3800 18440 3810
rect 18360 3790 18440 3800
rect 18500 3740 18580 3750
rect 18500 3730 18510 3740
rect 18360 3680 18510 3730
rect 18500 3670 18510 3680
rect 18570 3670 18580 3740
rect 18500 3660 18580 3670
rect 18360 3610 18440 3620
rect 18360 3540 18370 3610
rect 18430 3600 18440 3610
rect 18430 3550 18580 3600
rect 18430 3540 18440 3550
rect 18360 3530 18440 3540
rect 18500 3480 18580 3490
rect 18500 3472 18510 3480
rect 18371 3470 18510 3472
rect 18360 3420 18510 3470
rect 18500 3410 18510 3420
rect 18570 3410 18580 3480
rect 18500 3400 18580 3410
rect 18360 3360 18440 3370
rect 18360 3290 18370 3360
rect 18430 3350 18440 3360
rect 18430 3300 18580 3350
rect 18430 3298 18571 3300
rect 18430 3290 18440 3298
rect 18360 3280 18440 3290
rect 18500 3230 18580 3240
rect 18500 3220 18510 3230
rect 18360 3170 18510 3220
rect 18500 3160 18510 3170
rect 18570 3160 18580 3230
rect 18500 3150 18580 3160
rect 18360 3100 18440 3110
rect 18360 3030 18370 3100
rect 18430 3090 18440 3100
rect 18430 3040 18580 3090
rect 18430 3030 18440 3040
rect 18360 3020 18440 3030
rect 18500 2970 18580 2980
rect 18500 2960 18510 2970
rect 18360 2910 18510 2960
rect 18500 2900 18510 2910
rect 18570 2900 18580 2970
rect 18500 2890 18580 2900
rect 18360 2840 18440 2850
rect 18360 2770 18370 2840
rect 18430 2832 18440 2840
rect 18430 2830 18571 2832
rect 18430 2780 18580 2830
rect 18430 2770 18440 2780
rect 18360 2760 18440 2770
rect 18500 2720 18580 2730
rect 18500 2710 18510 2720
rect 18360 2650 18510 2710
rect 18570 2650 18580 2720
rect 18500 2640 18580 2650
rect 18360 2590 18440 2600
rect 18360 2520 18370 2590
rect 18430 2580 18440 2590
rect 18430 2530 18580 2580
rect 18430 2520 18440 2530
rect 18360 2510 18440 2520
rect 18500 2460 18580 2470
rect 18500 2450 18510 2460
rect 18360 2400 18510 2450
rect 18500 2390 18510 2400
rect 18570 2390 18580 2460
rect 18500 2380 18580 2390
rect 18360 2330 18440 2340
rect 18360 2260 18370 2330
rect 18430 2320 18440 2330
rect 18430 2270 18580 2320
rect 18430 2260 18440 2270
rect 18360 2250 18440 2260
rect 18500 2200 18580 2210
rect 18360 2140 18510 2200
rect 18500 2130 18510 2140
rect 18570 2130 18580 2200
rect 18500 2120 18580 2130
rect 18360 2080 18440 2090
rect 18360 2010 18370 2080
rect 18430 2070 18440 2080
rect 18430 2010 18580 2070
rect 18360 2000 18440 2010
rect 18500 1950 18580 1960
rect 18500 1940 18510 1950
rect 18360 1890 18510 1940
rect 18500 1880 18510 1890
rect 18570 1880 18580 1950
rect 18500 1870 18580 1880
rect 18360 1820 18440 1830
rect 18360 1750 18370 1820
rect 18430 1810 18440 1820
rect 18430 1760 18580 1810
rect 18430 1750 18440 1760
rect 18360 1740 18440 1750
rect 18500 1690 18580 1700
rect 18500 1680 18510 1690
rect 18360 1630 18510 1680
rect 18500 1620 18510 1630
rect 18570 1620 18580 1690
rect 18500 1610 18580 1620
rect 18360 1560 18440 1570
rect 18360 1490 18370 1560
rect 18430 1552 18440 1560
rect 18430 1550 18571 1552
rect 18430 1510 18580 1550
rect 18430 1506 18571 1510
rect 18430 1490 18440 1506
rect 18360 1480 18440 1490
rect 18500 1430 18580 1440
rect 18360 1380 18510 1430
rect 18371 1378 18510 1380
rect 18500 1360 18510 1378
rect 18570 1360 18580 1430
rect 18500 1350 18580 1360
rect 18360 1310 18440 1320
rect 18360 1240 18370 1310
rect 18430 1300 18440 1310
rect 18610 1310 18670 4310
rect 19200 2215 19770 4790
rect 19200 1840 19235 2215
rect 19725 1840 19770 2215
rect 20070 1845 20130 6160
rect 20160 6120 20250 6130
rect 20160 6060 20170 6120
rect 20240 6110 20250 6120
rect 20240 6070 20380 6110
rect 20240 6060 20250 6070
rect 20160 6050 20250 6060
rect 20290 5990 20380 6000
rect 20290 5980 20300 5990
rect 20160 5940 20300 5980
rect 20290 5930 20300 5940
rect 20370 5930 20380 5990
rect 20290 5920 20380 5930
rect 20160 5860 20250 5870
rect 20160 5800 20170 5860
rect 20240 5850 20250 5860
rect 20240 5810 20380 5850
rect 20240 5800 20250 5810
rect 20160 5790 20250 5800
rect 20290 5730 20380 5740
rect 20290 5720 20300 5730
rect 20160 5680 20300 5720
rect 20290 5670 20300 5680
rect 20370 5670 20380 5730
rect 20290 5660 20380 5670
rect 20160 5610 20250 5620
rect 20160 5550 20170 5610
rect 20240 5600 20250 5610
rect 20240 5550 20380 5600
rect 20160 5540 20250 5550
rect 20290 5480 20380 5490
rect 20290 5470 20300 5480
rect 20160 5420 20300 5470
rect 20370 5420 20380 5480
rect 20290 5410 20380 5420
rect 20160 5350 20250 5360
rect 20160 5290 20170 5350
rect 20240 5340 20250 5350
rect 20240 5300 20380 5340
rect 20240 5290 20250 5300
rect 20160 5280 20250 5290
rect 20290 5220 20380 5230
rect 20290 5210 20300 5220
rect 20160 5170 20300 5210
rect 20290 5160 20300 5170
rect 20370 5160 20380 5220
rect 20290 5150 20380 5160
rect 20160 5090 20250 5100
rect 20160 5030 20170 5090
rect 20240 5040 20380 5090
rect 20240 5030 20250 5040
rect 20160 5020 20250 5030
rect 20290 4960 20380 4970
rect 20160 4910 20300 4960
rect 20290 4900 20300 4910
rect 20370 4900 20380 4960
rect 20290 4890 20380 4900
rect 20160 4830 20250 4840
rect 20160 4770 20170 4830
rect 20240 4780 20380 4830
rect 20240 4770 20250 4780
rect 20160 4760 20250 4770
rect 20290 4710 20380 4720
rect 20290 4700 20300 4710
rect 20160 4660 20300 4700
rect 20290 4650 20300 4660
rect 20370 4650 20380 4710
rect 20290 4640 20380 4650
rect 20160 4580 20250 4590
rect 20160 4520 20170 4580
rect 20240 4570 20250 4580
rect 20240 4530 20380 4570
rect 20240 4520 20250 4530
rect 20160 4510 20250 4520
rect 20290 4450 20380 4460
rect 20290 4440 20300 4450
rect 20160 4400 20300 4440
rect 20290 4390 20300 4400
rect 20370 4390 20380 4450
rect 20290 4380 20380 4390
rect 20160 4320 20250 4330
rect 20160 4260 20170 4320
rect 20240 4270 20380 4320
rect 20240 4260 20250 4270
rect 20160 4250 20250 4260
rect 20290 4200 20380 4210
rect 20290 4190 20300 4200
rect 20160 4140 20300 4190
rect 20370 4140 20380 4200
rect 20290 4130 20380 4140
rect 20290 3865 20380 3875
rect 20160 3815 20300 3865
rect 20290 3805 20300 3815
rect 20370 3805 20380 3865
rect 20290 3795 20380 3805
rect 20160 3745 20250 3755
rect 20160 3685 20170 3745
rect 20240 3735 20250 3745
rect 20240 3685 20380 3735
rect 20160 3675 20250 3685
rect 20290 3615 20380 3625
rect 20290 3605 20300 3615
rect 20160 3565 20300 3605
rect 20169 3559 20300 3565
rect 20290 3555 20300 3559
rect 20370 3555 20380 3615
rect 20290 3545 20380 3555
rect 20160 3485 20250 3495
rect 20160 3425 20170 3485
rect 20240 3477 20250 3485
rect 20240 3475 20369 3477
rect 20240 3435 20380 3475
rect 20240 3431 20369 3435
rect 20240 3425 20250 3431
rect 20160 3415 20250 3425
rect 20290 3355 20380 3365
rect 20290 3349 20300 3355
rect 20169 3345 20300 3349
rect 20160 3305 20300 3345
rect 20169 3303 20300 3305
rect 20290 3295 20300 3303
rect 20370 3295 20380 3355
rect 20290 3285 20380 3295
rect 20160 3235 20250 3245
rect 20160 3175 20170 3235
rect 20240 3225 20250 3235
rect 20240 3175 20380 3225
rect 20160 3165 20250 3175
rect 20290 3105 20380 3115
rect 20290 3095 20300 3105
rect 20160 3045 20300 3095
rect 20370 3045 20380 3105
rect 20290 3035 20380 3045
rect 20160 2975 20250 2985
rect 20160 2915 20170 2975
rect 20240 2965 20250 2975
rect 20240 2915 20380 2965
rect 20160 2905 20250 2915
rect 20290 2845 20380 2855
rect 20290 2837 20300 2845
rect 20169 2835 20300 2837
rect 20160 2795 20300 2835
rect 20169 2791 20300 2795
rect 20290 2785 20300 2791
rect 20370 2785 20380 2845
rect 20290 2775 20380 2785
rect 20160 2715 20250 2725
rect 20160 2655 20170 2715
rect 20240 2709 20250 2715
rect 20240 2705 20369 2709
rect 20240 2665 20380 2705
rect 20240 2663 20369 2665
rect 20240 2655 20250 2663
rect 20160 2645 20250 2655
rect 20290 2585 20380 2595
rect 20160 2535 20300 2585
rect 20290 2525 20300 2535
rect 20370 2525 20380 2585
rect 20290 2515 20380 2525
rect 20160 2455 20250 2465
rect 20160 2395 20170 2455
rect 20240 2405 20380 2455
rect 20240 2395 20250 2405
rect 20160 2385 20250 2395
rect 20290 2335 20380 2345
rect 20290 2325 20300 2335
rect 20160 2285 20300 2325
rect 20169 2279 20300 2285
rect 20290 2275 20300 2279
rect 20370 2275 20380 2335
rect 20290 2265 20380 2275
rect 20160 2205 20250 2215
rect 20160 2145 20170 2205
rect 20240 2197 20250 2205
rect 20240 2195 20369 2197
rect 20240 2155 20380 2195
rect 20240 2151 20369 2155
rect 20240 2145 20250 2151
rect 20160 2135 20250 2145
rect 20290 2075 20380 2085
rect 20290 2069 20300 2075
rect 20169 2065 20300 2069
rect 20160 2025 20300 2065
rect 20169 2023 20300 2025
rect 20290 2015 20300 2023
rect 20370 2015 20380 2075
rect 20290 2005 20380 2015
rect 20160 1945 20250 1955
rect 20160 1885 20170 1945
rect 20240 1941 20250 1945
rect 20240 1935 20369 1941
rect 20240 1895 20380 1935
rect 20240 1885 20250 1895
rect 20160 1875 20250 1885
rect 20410 1845 20470 6160
rect 20820 5520 21340 5580
rect 20820 4180 20880 5520
rect 20910 5480 21000 5490
rect 20910 5420 20920 5480
rect 20990 5470 21000 5480
rect 20990 5420 21130 5470
rect 20910 5410 21000 5420
rect 21040 5350 21130 5360
rect 21040 5340 21050 5350
rect 20910 5290 21050 5340
rect 21120 5290 21130 5350
rect 21040 5280 21130 5290
rect 20910 5220 21000 5230
rect 20910 5160 20920 5220
rect 20990 5170 21130 5220
rect 20990 5160 21000 5170
rect 20910 5150 21000 5160
rect 21040 5100 21130 5110
rect 21040 5090 21050 5100
rect 20910 5040 21050 5090
rect 21040 5030 21050 5040
rect 21120 5030 21130 5100
rect 21040 5020 21130 5030
rect 20910 4970 21000 4980
rect 20910 4910 20920 4970
rect 20990 4960 21000 4970
rect 20990 4910 21130 4960
rect 20910 4900 21000 4910
rect 21040 4840 21130 4850
rect 21040 4830 21050 4840
rect 20910 4780 21050 4830
rect 21120 4780 21130 4840
rect 21040 4770 21130 4780
rect 20910 4710 21000 4720
rect 20910 4650 20920 4710
rect 20990 4700 21000 4710
rect 20990 4660 21130 4700
rect 20990 4650 21000 4660
rect 20910 4640 21000 4650
rect 21040 4580 21130 4590
rect 21040 4570 21050 4580
rect 20910 4530 21050 4570
rect 21040 4520 21050 4530
rect 21120 4520 21130 4580
rect 21040 4510 21130 4520
rect 20910 4450 21000 4460
rect 20910 4390 20920 4450
rect 20990 4400 21130 4450
rect 20990 4390 21000 4400
rect 20910 4380 21000 4390
rect 21040 4320 21130 4330
rect 20910 4270 21050 4320
rect 21040 4260 21050 4270
rect 21120 4260 21130 4320
rect 21040 4250 21130 4260
rect 20910 4200 21000 4210
rect 20910 4140 20920 4200
rect 20990 4190 21000 4200
rect 20990 4140 21130 4190
rect 21160 4180 21220 5520
rect 20910 4130 21000 4140
rect 20910 3875 21000 3885
rect 20820 2495 20880 3835
rect 20910 3815 20920 3875
rect 20990 3825 21130 3875
rect 20990 3815 21000 3825
rect 20910 3805 21000 3815
rect 21040 3755 21130 3765
rect 21040 3745 21050 3755
rect 20910 3695 21050 3745
rect 21120 3695 21130 3755
rect 21040 3685 21130 3695
rect 20910 3625 21000 3635
rect 20910 3565 20920 3625
rect 20990 3615 21000 3625
rect 20990 3565 21130 3615
rect 20910 3555 21000 3565
rect 21040 3495 21130 3505
rect 21040 3487 21050 3495
rect 20919 3485 21050 3487
rect 20910 3445 21050 3485
rect 20919 3441 21050 3445
rect 21040 3435 21050 3441
rect 21120 3435 21130 3495
rect 21040 3425 21130 3435
rect 20910 3365 21000 3375
rect 20910 3305 20920 3365
rect 20990 3359 21000 3365
rect 20990 3355 21119 3359
rect 20990 3315 21130 3355
rect 20990 3313 21119 3315
rect 20990 3305 21000 3313
rect 20910 3295 21000 3305
rect 21040 3235 21130 3245
rect 20910 3185 21050 3235
rect 21040 3175 21050 3185
rect 21120 3175 21130 3235
rect 21040 3165 21130 3175
rect 20910 3105 21000 3115
rect 20910 3045 20920 3105
rect 20990 3055 21130 3105
rect 20990 3045 21000 3055
rect 20910 3035 21000 3045
rect 21040 2985 21130 2995
rect 21040 2975 21050 2985
rect 20910 2925 21050 2975
rect 21040 2915 21050 2925
rect 21120 2915 21130 2985
rect 21040 2905 21130 2915
rect 20910 2855 21000 2865
rect 20910 2795 20920 2855
rect 20990 2847 21000 2855
rect 20990 2845 21119 2847
rect 20990 2795 21130 2845
rect 20910 2785 21000 2795
rect 21040 2725 21130 2735
rect 20910 2675 21050 2725
rect 20919 2673 21050 2675
rect 21040 2665 21050 2673
rect 21120 2665 21130 2725
rect 21040 2655 21130 2665
rect 20910 2595 21000 2605
rect 20910 2535 20920 2595
rect 20990 2545 21130 2595
rect 20990 2535 21000 2545
rect 20910 2525 21000 2535
rect 21160 2495 21220 3835
rect 20820 2435 21340 2495
rect 19200 1800 19770 1840
rect 18430 1250 18580 1300
rect 18430 1240 18440 1250
rect 18360 1230 18440 1240
rect 18500 1180 18580 1190
rect 18500 1170 18510 1180
rect 18360 1120 18510 1170
rect 18500 1110 18510 1120
rect 18570 1110 18580 1180
rect 18500 1100 18580 1110
rect 18360 1050 18440 1060
rect 18360 980 18370 1050
rect 18430 1040 18440 1050
rect 18430 990 18580 1040
rect 18430 980 18440 990
rect 18360 970 18440 980
rect 18500 920 18580 930
rect 18500 912 18510 920
rect 18371 910 18510 912
rect 18360 860 18510 910
rect 18500 850 18510 860
rect 18570 850 18580 920
rect 18500 840 18580 850
rect 18610 880 19240 1310
rect 18360 800 18440 810
rect 18360 730 18370 800
rect 18430 790 18440 800
rect 18430 730 18580 790
rect 18360 720 18440 730
rect 18500 670 18580 680
rect 18500 660 18510 670
rect 18360 610 18510 660
rect 18500 600 18510 610
rect 18570 600 18580 670
rect 18500 590 18580 600
rect 18360 540 18440 550
rect 18360 470 18370 540
rect 18430 530 18440 540
rect 18430 480 18580 530
rect 18430 470 18440 480
rect 18360 460 18440 470
rect 18500 410 18580 420
rect 18500 400 18510 410
rect 17780 350 17930 400
rect 18360 350 18510 400
rect 17780 340 17790 350
rect 17710 330 17790 340
rect 18500 340 18510 350
rect 18570 340 18580 410
rect 18610 400 18670 880
rect 18500 330 18580 340
rect 17390 -130 17495 -125
rect 17390 -160 17400 -130
rect 16985 -185 17400 -160
rect 17480 -160 17495 -130
rect 17775 -135 17880 -120
rect 17775 -160 17785 -135
rect 17480 -185 17785 -160
rect 16985 -190 17785 -185
rect 17865 -160 17880 -135
rect 17980 -130 18085 -120
rect 17980 -160 17995 -130
rect 17865 -185 17995 -160
rect 18075 -160 18085 -130
rect 18075 -185 19305 -160
rect 17865 -190 19305 -185
rect 16985 -210 19305 -190
rect 16985 -365 17040 -240
rect 17070 -250 17145 -240
rect 17070 -305 17080 -250
rect 17135 -305 17145 -250
rect 17070 -315 17145 -305
rect 16970 -375 17045 -365
rect 16970 -430 16980 -375
rect 17035 -430 17045 -375
rect 16970 -440 17045 -430
rect 17080 -440 17135 -315
rect 17175 -365 17230 -240
rect 17260 -250 17335 -240
rect 17260 -305 17270 -250
rect 17325 -305 17335 -250
rect 17260 -315 17335 -305
rect 17165 -375 17240 -365
rect 17165 -430 17175 -375
rect 17230 -430 17240 -375
rect 17165 -440 17240 -430
rect 17275 -440 17325 -315
rect 17370 -365 17425 -240
rect 17455 -250 17530 -240
rect 17455 -305 17465 -250
rect 17520 -305 17530 -250
rect 17455 -315 17530 -305
rect 17360 -375 17435 -365
rect 17360 -430 17370 -375
rect 17425 -430 17435 -375
rect 17360 -440 17435 -430
rect 17465 -440 17520 -315
rect 17560 -365 17615 -240
rect 17645 -250 17720 -240
rect 17645 -305 17655 -250
rect 17710 -305 17720 -250
rect 17645 -315 17720 -305
rect 17550 -375 17625 -365
rect 17550 -430 17560 -375
rect 17615 -430 17625 -375
rect 17550 -440 17625 -430
rect 17655 -440 17710 -315
rect 17755 -365 17810 -240
rect 17840 -250 17915 -240
rect 17840 -305 17850 -250
rect 17905 -305 17915 -250
rect 17840 -315 17915 -305
rect 17740 -375 17815 -365
rect 17740 -430 17750 -375
rect 17805 -430 17815 -375
rect 17740 -440 17815 -430
rect 17850 -440 17905 -315
rect 17945 -365 18000 -240
rect 17935 -375 18010 -365
rect 17935 -430 17945 -375
rect 18000 -430 18010 -375
rect 17935 -440 18010 -430
rect 18125 -470 18165 -210
rect 18290 -365 18345 -240
rect 18375 -250 18450 -240
rect 18375 -305 18385 -250
rect 18440 -305 18450 -250
rect 18375 -315 18450 -305
rect 18280 -375 18355 -365
rect 18280 -430 18290 -375
rect 18345 -430 18355 -375
rect 18280 -440 18355 -430
rect 18385 -440 18440 -315
rect 18480 -365 18535 -240
rect 18570 -250 18645 -240
rect 18570 -305 18580 -250
rect 18635 -305 18645 -250
rect 18570 -315 18645 -305
rect 18475 -375 18550 -365
rect 18475 -430 18485 -375
rect 18540 -430 18550 -375
rect 18475 -440 18550 -430
rect 18580 -440 18635 -315
rect 18675 -365 18730 -240
rect 18760 -250 18835 -240
rect 18760 -305 18770 -250
rect 18825 -305 18835 -250
rect 18760 -315 18835 -305
rect 18665 -375 18740 -365
rect 18665 -430 18675 -375
rect 18730 -430 18740 -375
rect 18665 -440 18740 -430
rect 18770 -440 18825 -315
rect 18865 -365 18920 -240
rect 18955 -250 19030 -240
rect 18955 -305 18965 -250
rect 19020 -305 19030 -250
rect 18955 -315 19030 -305
rect 18855 -375 18930 -365
rect 18855 -430 18865 -375
rect 18920 -430 18930 -375
rect 18855 -440 18930 -430
rect 18965 -440 19015 -315
rect 19060 -365 19115 -240
rect 19145 -250 19220 -240
rect 19145 -305 19155 -250
rect 19210 -305 19220 -250
rect 19145 -315 19220 -305
rect 19050 -375 19125 -365
rect 19050 -430 19060 -375
rect 19115 -430 19125 -375
rect 19050 -440 19125 -430
rect 19155 -440 19210 -315
rect 19250 -365 19305 -240
rect 19245 -375 19320 -365
rect 19245 -430 19255 -375
rect 19310 -430 19320 -375
rect 19245 -440 19320 -430
rect 16980 -520 19310 -470
<< via1 >>
rect 17320 7050 17390 7110
rect 17450 6920 17520 6980
rect 17320 6790 17390 6850
rect 17450 6660 17520 6720
rect 17320 6530 17390 6590
rect 17450 6400 17520 6460
rect 17320 6270 17390 6330
rect 17450 6150 17520 6210
rect 17320 6020 17390 6080
rect 17450 5900 17520 5960
rect 17320 5770 17390 5830
rect 17450 5640 17520 5700
rect 17320 5510 17390 5570
rect 17450 5380 17520 5440
rect 17320 5250 17390 5310
rect 17970 7050 18040 7110
rect 18100 6920 18170 6980
rect 17970 6790 18040 6850
rect 18100 6660 18170 6720
rect 17970 6530 18040 6590
rect 18100 6400 18170 6460
rect 17970 6270 18040 6330
rect 18100 6150 18170 6210
rect 17970 6020 18040 6080
rect 18100 5900 18170 5960
rect 17970 5770 18040 5830
rect 18100 5640 18170 5700
rect 17970 5510 18040 5570
rect 18100 5380 18170 5440
rect 17970 5250 18040 5310
rect 18620 7050 18690 7110
rect 18750 6920 18820 6980
rect 18620 6790 18690 6850
rect 18750 6660 18820 6720
rect 18620 6530 18690 6590
rect 18750 6400 18820 6460
rect 18620 6270 18690 6330
rect 18750 6150 18820 6210
rect 18620 6020 18690 6080
rect 18750 5900 18820 5960
rect 18620 5770 18690 5830
rect 18750 5640 18820 5700
rect 18620 5510 18690 5570
rect 18750 5380 18820 5440
rect 18620 5250 18690 5310
rect 19235 6325 19740 6710
rect 17450 5120 17520 5180
rect 18100 5120 18170 5180
rect 18750 5120 18820 5180
rect 17720 4180 17780 4250
rect 17860 4050 17920 4120
rect 17720 3920 17780 3990
rect 17860 3800 17920 3870
rect 17720 3670 17780 3740
rect 17860 3540 17920 3610
rect 17720 3410 17780 3480
rect 17860 3290 17920 3360
rect 17720 3160 17780 3230
rect 17860 3030 17920 3100
rect 17720 2900 17780 2970
rect 17860 2770 17920 2840
rect 17720 2650 17780 2720
rect 17860 2520 17920 2590
rect 17720 2390 17780 2460
rect 17860 2260 17920 2330
rect 17720 2130 17780 2200
rect 17860 2010 17920 2080
rect 17720 1880 17780 1950
rect 17860 1750 17920 1820
rect 17720 1620 17780 1690
rect 17860 1490 17920 1560
rect 17720 1360 17780 1430
rect 17860 1240 17920 1310
rect 17720 1110 17780 1180
rect 17860 980 17920 1050
rect 17720 850 17780 920
rect 17860 730 17920 800
rect 17720 600 17780 670
rect 17860 470 17920 540
rect 17720 340 17780 410
rect 18510 4180 18570 4250
rect 18370 4050 18430 4120
rect 18510 3920 18570 3990
rect 18370 3800 18430 3870
rect 18510 3670 18570 3740
rect 18370 3540 18430 3610
rect 18510 3410 18570 3480
rect 18370 3290 18430 3360
rect 18510 3160 18570 3230
rect 18370 3030 18430 3100
rect 18510 2900 18570 2970
rect 18370 2770 18430 2840
rect 18510 2650 18570 2720
rect 18370 2520 18430 2590
rect 18510 2390 18570 2460
rect 18370 2260 18430 2330
rect 18510 2130 18570 2200
rect 18370 2010 18430 2080
rect 18510 1880 18570 1950
rect 18370 1750 18430 1820
rect 18510 1620 18570 1690
rect 18370 1490 18430 1560
rect 18510 1360 18570 1430
rect 18370 1240 18430 1310
rect 19235 1840 19725 2215
rect 20170 6060 20240 6120
rect 20300 5930 20370 5990
rect 20170 5800 20240 5860
rect 20300 5670 20370 5730
rect 20170 5550 20240 5610
rect 20300 5420 20370 5480
rect 20170 5290 20240 5350
rect 20300 5160 20370 5220
rect 20170 5030 20240 5090
rect 20300 4900 20370 4960
rect 20170 4770 20240 4830
rect 20300 4650 20370 4710
rect 20170 4520 20240 4580
rect 20300 4390 20370 4450
rect 20170 4260 20240 4320
rect 20300 4140 20370 4200
rect 20300 3805 20370 3865
rect 20170 3685 20240 3745
rect 20300 3555 20370 3615
rect 20170 3425 20240 3485
rect 20300 3295 20370 3355
rect 20170 3175 20240 3235
rect 20300 3045 20370 3105
rect 20170 2915 20240 2975
rect 20300 2785 20370 2845
rect 20170 2655 20240 2715
rect 20300 2525 20370 2585
rect 20170 2395 20240 2455
rect 20300 2275 20370 2335
rect 20170 2145 20240 2205
rect 20300 2015 20370 2075
rect 20170 1885 20240 1945
rect 20920 5420 20990 5480
rect 21050 5290 21120 5350
rect 20920 5160 20990 5220
rect 21050 5030 21120 5100
rect 20920 4910 20990 4970
rect 21050 4780 21120 4840
rect 20920 4650 20990 4710
rect 21050 4520 21120 4580
rect 20920 4390 20990 4450
rect 21050 4260 21120 4320
rect 20920 4140 20990 4200
rect 20920 3815 20990 3875
rect 21050 3695 21120 3755
rect 20920 3565 20990 3625
rect 21050 3435 21120 3495
rect 20920 3305 20990 3365
rect 21050 3175 21120 3235
rect 20920 3045 20990 3105
rect 21050 2915 21120 2985
rect 20920 2795 20990 2855
rect 21050 2665 21120 2725
rect 20920 2535 20990 2595
rect 18510 1110 18570 1180
rect 18370 980 18430 1050
rect 18510 850 18570 920
rect 19240 910 19750 1280
rect 18370 730 18430 800
rect 18510 600 18570 670
rect 18370 470 18430 540
rect 18510 340 18570 410
rect 17400 -185 17480 -130
rect 17785 -190 17865 -135
rect 17995 -185 18075 -130
rect 17080 -305 17135 -250
rect 16980 -430 17035 -375
rect 17270 -305 17325 -250
rect 17175 -430 17230 -375
rect 17465 -305 17520 -250
rect 17370 -430 17425 -375
rect 17655 -305 17710 -250
rect 17560 -430 17615 -375
rect 17850 -305 17905 -250
rect 17750 -430 17805 -375
rect 17945 -430 18000 -375
rect 18385 -305 18440 -250
rect 18290 -430 18345 -375
rect 18580 -305 18635 -250
rect 18485 -430 18540 -375
rect 18770 -305 18825 -250
rect 18675 -430 18730 -375
rect 18965 -305 19020 -250
rect 18865 -430 18920 -375
rect 19155 -305 19210 -250
rect 19060 -430 19115 -375
rect 19255 -430 19310 -375
<< metal2 >>
rect 17440 7265 17720 7275
rect 17440 7150 17450 7265
rect 17705 7150 17720 7265
rect 17100 7110 17400 7120
rect 17100 7050 17320 7110
rect 17390 7050 17400 7110
rect 17100 6850 17400 7050
rect 17100 6790 17320 6850
rect 17390 6790 17400 6850
rect 17100 6590 17400 6790
rect 17100 6530 17320 6590
rect 17390 6530 17400 6590
rect 17100 6330 17400 6530
rect 17100 6270 17320 6330
rect 17390 6270 17400 6330
rect 17100 6080 17400 6270
rect 17100 6020 17320 6080
rect 17390 6020 17400 6080
rect 17100 5830 17400 6020
rect 17100 5770 17320 5830
rect 17390 5770 17400 5830
rect 17100 5570 17400 5770
rect 17100 5510 17320 5570
rect 17390 5510 17400 5570
rect 17100 5310 17400 5510
rect 17100 5250 17320 5310
rect 17390 5250 17400 5310
rect 17100 5000 17400 5250
rect 17440 6980 17720 7150
rect 18090 7265 18370 7275
rect 18090 7150 18105 7265
rect 18360 7150 18370 7265
rect 17440 6920 17450 6980
rect 17520 6920 17720 6980
rect 17440 6720 17720 6920
rect 17440 6660 17450 6720
rect 17520 6660 17720 6720
rect 17440 6460 17720 6660
rect 17440 6400 17450 6460
rect 17520 6400 17720 6460
rect 17440 6210 17720 6400
rect 17440 6150 17450 6210
rect 17520 6150 17720 6210
rect 17440 5960 17720 6150
rect 17440 5900 17450 5960
rect 17520 5900 17720 5960
rect 17440 5700 17720 5900
rect 17440 5640 17450 5700
rect 17520 5640 17720 5700
rect 17440 5440 17720 5640
rect 17440 5380 17450 5440
rect 17520 5380 17720 5440
rect 17440 5180 17720 5380
rect 17440 5120 17450 5180
rect 17520 5120 17720 5180
rect 17440 5110 17720 5120
rect 17760 7110 18050 7120
rect 17760 7050 17970 7110
rect 18040 7050 18050 7110
rect 17760 6850 18050 7050
rect 17760 6790 17970 6850
rect 18040 6790 18050 6850
rect 17760 6590 18050 6790
rect 17760 6530 17970 6590
rect 18040 6530 18050 6590
rect 17760 6330 18050 6530
rect 17760 6270 17970 6330
rect 18040 6270 18050 6330
rect 17760 6080 18050 6270
rect 17760 6020 17970 6080
rect 18040 6020 18050 6080
rect 17760 5830 18050 6020
rect 17760 5770 17970 5830
rect 18040 5770 18050 5830
rect 17760 5570 18050 5770
rect 17760 5510 17970 5570
rect 18040 5510 18050 5570
rect 17760 5310 18050 5510
rect 17760 5250 17970 5310
rect 18040 5250 18050 5310
rect 17760 5000 18050 5250
rect 18090 6980 18370 7150
rect 18740 7265 19020 7275
rect 18740 7150 18750 7265
rect 19005 7150 19020 7265
rect 18090 6920 18100 6980
rect 18170 6920 18370 6980
rect 18090 6720 18370 6920
rect 18090 6660 18100 6720
rect 18170 6660 18370 6720
rect 18090 6460 18370 6660
rect 18090 6400 18100 6460
rect 18170 6400 18370 6460
rect 18090 6210 18370 6400
rect 18090 6150 18100 6210
rect 18170 6150 18370 6210
rect 18090 5960 18370 6150
rect 18090 5900 18100 5960
rect 18170 5900 18370 5960
rect 18090 5700 18370 5900
rect 18090 5640 18100 5700
rect 18170 5640 18370 5700
rect 18090 5440 18370 5640
rect 18090 5380 18100 5440
rect 18170 5380 18370 5440
rect 18090 5180 18370 5380
rect 18090 5120 18100 5180
rect 18170 5120 18370 5180
rect 18090 5110 18370 5120
rect 18410 7110 18700 7120
rect 18410 7050 18620 7110
rect 18690 7050 18700 7110
rect 18410 6850 18700 7050
rect 18410 6790 18620 6850
rect 18690 6790 18700 6850
rect 18410 6590 18700 6790
rect 18410 6530 18620 6590
rect 18690 6530 18700 6590
rect 18410 6330 18700 6530
rect 18410 6270 18620 6330
rect 18690 6270 18700 6330
rect 18410 6080 18700 6270
rect 18410 6020 18620 6080
rect 18690 6020 18700 6080
rect 18410 5830 18700 6020
rect 18410 5770 18620 5830
rect 18690 5770 18700 5830
rect 18410 5570 18700 5770
rect 18410 5510 18620 5570
rect 18690 5510 18700 5570
rect 18410 5310 18700 5510
rect 18410 5250 18620 5310
rect 18690 5250 18700 5310
rect 18410 5000 18700 5250
rect 18740 6980 19020 7150
rect 18740 6920 18750 6980
rect 18820 6920 19020 6980
rect 18740 6720 19020 6920
rect 18740 6660 18750 6720
rect 18820 6660 19020 6720
rect 18740 6460 19020 6660
rect 18740 6400 18750 6460
rect 18820 6400 19020 6460
rect 18740 6210 19020 6400
rect 19210 6710 21340 6745
rect 19210 6325 19235 6710
rect 19740 6325 21340 6710
rect 19210 6300 21340 6325
rect 18740 6150 18750 6210
rect 18820 6150 19020 6210
rect 18740 5960 19020 6150
rect 18740 5900 18750 5960
rect 18820 5900 19020 5960
rect 18740 5700 19020 5900
rect 18740 5640 18750 5700
rect 18820 5640 19020 5700
rect 18740 5440 19020 5640
rect 18740 5380 18750 5440
rect 18820 5380 19020 5440
rect 18740 5180 19020 5380
rect 18740 5120 18750 5180
rect 18820 5120 19020 5180
rect 18740 5110 19020 5120
rect 19950 6135 20250 6150
rect 19950 5925 19970 6135
rect 20230 6120 20250 6135
rect 20240 6060 20250 6120
rect 20230 5925 20250 6060
rect 19950 5860 20250 5925
rect 19950 5800 20170 5860
rect 20240 5800 20250 5860
rect 19950 5610 20250 5800
rect 19950 5550 20170 5610
rect 20240 5550 20250 5610
rect 19950 5350 20250 5550
rect 19950 5290 20170 5350
rect 20240 5290 20250 5350
rect 17100 4400 18700 5000
rect 19950 5090 20250 5290
rect 19950 5030 20170 5090
rect 20240 5030 20250 5090
rect 19950 4830 20250 5030
rect 19950 4770 20170 4830
rect 20240 4770 20250 4830
rect 19950 4580 20250 4770
rect 19950 4520 20170 4580
rect 20240 4520 20250 4580
rect 17190 4250 17790 4260
rect 17190 4180 17720 4250
rect 17780 4180 17790 4250
rect 17190 3990 17790 4180
rect 17190 3920 17720 3990
rect 17780 3920 17790 3990
rect 17190 3740 17790 3920
rect 17190 3670 17720 3740
rect 17780 3670 17790 3740
rect 17190 3480 17790 3670
rect 17190 3410 17720 3480
rect 17780 3410 17790 3480
rect 17190 3230 17790 3410
rect 17190 3160 17720 3230
rect 17780 3160 17790 3230
rect 17190 2970 17790 3160
rect 17190 2900 17720 2970
rect 17780 2900 17790 2970
rect 17190 2720 17790 2900
rect 17190 2650 17720 2720
rect 17780 2650 17790 2720
rect 17190 2460 17790 2650
rect 17190 2390 17720 2460
rect 17780 2390 17790 2460
rect 17190 2200 17790 2390
rect 17190 2130 17720 2200
rect 17780 2130 17790 2200
rect 17190 1950 17790 2130
rect 17190 1880 17720 1950
rect 17780 1880 17790 1950
rect 17190 1690 17790 1880
rect 17190 1620 17720 1690
rect 17780 1620 17790 1690
rect 17190 1430 17790 1620
rect 17190 1360 17720 1430
rect 17780 1360 17790 1430
rect 17190 1180 17790 1360
rect 17190 1110 17720 1180
rect 17780 1110 17790 1180
rect 17190 920 17790 1110
rect 17190 850 17720 920
rect 17780 850 17790 920
rect 17190 670 17790 850
rect 17190 600 17720 670
rect 17780 600 17790 670
rect 17190 410 17790 600
rect 17850 4120 18440 4400
rect 19950 4320 20250 4520
rect 19950 4260 20170 4320
rect 20240 4260 20250 4320
rect 17850 4050 17860 4120
rect 17920 4050 18370 4120
rect 18430 4050 18440 4120
rect 17850 3870 18440 4050
rect 17850 3800 17860 3870
rect 17920 3800 18370 3870
rect 18430 3800 18440 3870
rect 17850 3610 18440 3800
rect 17850 3540 17860 3610
rect 17920 3540 18370 3610
rect 18430 3540 18440 3610
rect 17850 3360 18440 3540
rect 17850 3290 17860 3360
rect 17920 3290 18370 3360
rect 18430 3290 18440 3360
rect 17850 3100 18440 3290
rect 17850 3030 17860 3100
rect 17920 3030 18370 3100
rect 18430 3030 18440 3100
rect 17850 2840 18440 3030
rect 17850 2770 17860 2840
rect 17920 2770 18370 2840
rect 18430 2770 18440 2840
rect 17850 2590 18440 2770
rect 17850 2520 17860 2590
rect 17920 2520 18370 2590
rect 18430 2520 18440 2590
rect 17850 2330 18440 2520
rect 17850 2260 17860 2330
rect 17920 2260 18370 2330
rect 18430 2260 18440 2330
rect 17850 2080 18440 2260
rect 17850 2010 17860 2080
rect 17920 2010 18370 2080
rect 18430 2010 18440 2080
rect 17850 1820 18440 2010
rect 17850 1750 17860 1820
rect 17920 1750 18370 1820
rect 18430 1750 18440 1820
rect 17850 1560 18440 1750
rect 17850 1490 17860 1560
rect 17920 1490 18370 1560
rect 18430 1490 18440 1560
rect 17850 1310 18440 1490
rect 17850 1240 17860 1310
rect 17920 1240 18370 1310
rect 18430 1240 18440 1310
rect 17850 1050 18440 1240
rect 17850 980 17860 1050
rect 17920 980 18370 1050
rect 18430 980 18440 1050
rect 17850 800 18440 980
rect 17850 730 17860 800
rect 17920 730 18370 800
rect 18430 730 18440 800
rect 17850 540 18440 730
rect 17850 470 17860 540
rect 17920 470 18370 540
rect 18430 470 18440 540
rect 17850 460 18440 470
rect 18500 4250 19100 4260
rect 18500 4180 18510 4250
rect 18570 4180 19100 4250
rect 18500 3990 19100 4180
rect 18500 3920 18510 3990
rect 18570 3920 19100 3990
rect 18500 3740 19100 3920
rect 18500 3670 18510 3740
rect 18570 3670 19100 3740
rect 18500 3480 19100 3670
rect 18500 3410 18510 3480
rect 18570 3410 19100 3480
rect 18500 3230 19100 3410
rect 18500 3160 18510 3230
rect 18570 3160 19100 3230
rect 18500 2970 19100 3160
rect 18500 2900 18510 2970
rect 18570 2900 19100 2970
rect 18500 2720 19100 2900
rect 18500 2650 18510 2720
rect 18570 2650 19100 2720
rect 18500 2460 19100 2650
rect 18500 2390 18510 2460
rect 18570 2390 19100 2460
rect 18500 2200 19100 2390
rect 19950 3745 20250 4260
rect 19950 3685 20170 3745
rect 20240 3685 20250 3745
rect 19950 3485 20250 3685
rect 19950 3425 20170 3485
rect 20240 3425 20250 3485
rect 19950 3235 20250 3425
rect 19950 3175 20170 3235
rect 20240 3175 20250 3235
rect 19950 2975 20250 3175
rect 19950 2915 20170 2975
rect 20240 2915 20250 2975
rect 19950 2715 20250 2915
rect 19950 2655 20170 2715
rect 20240 2655 20250 2715
rect 19950 2455 20250 2655
rect 19950 2395 20170 2455
rect 20240 2395 20250 2455
rect 18500 2130 18510 2200
rect 18570 2130 19100 2200
rect 18500 1950 19100 2130
rect 18500 1880 18510 1950
rect 18570 1880 19100 1950
rect 18500 1690 19100 1880
rect 19200 2215 19770 2255
rect 19200 1840 19235 2215
rect 19725 1840 19770 2215
rect 19950 2205 20250 2395
rect 19950 2145 20170 2205
rect 20240 2145 20250 2205
rect 19950 1945 20250 2145
rect 19950 1885 20170 1945
rect 20240 1885 20250 1945
rect 19950 1855 20250 1885
rect 20290 5990 20590 6150
rect 20290 5930 20300 5990
rect 20370 5930 20590 5990
rect 20290 5730 20590 5930
rect 20290 5670 20300 5730
rect 20370 5670 20590 5730
rect 20290 5480 20590 5670
rect 20290 5420 20300 5480
rect 20370 5420 20590 5480
rect 20290 5220 20590 5420
rect 20290 5160 20300 5220
rect 20370 5160 20590 5220
rect 20290 4960 20590 5160
rect 20290 4900 20300 4960
rect 20370 4900 20590 4960
rect 20290 4710 20590 4900
rect 20290 4650 20300 4710
rect 20370 4650 20590 4710
rect 20290 4450 20590 4650
rect 20290 4390 20300 4450
rect 20370 4390 20590 4450
rect 20290 4200 20590 4390
rect 20290 4140 20300 4200
rect 20370 4160 20590 4200
rect 20700 5480 21000 5490
rect 20700 5420 20920 5480
rect 20990 5420 21000 5480
rect 20700 5220 21000 5420
rect 20700 5160 20920 5220
rect 20990 5160 21000 5220
rect 20700 4970 21000 5160
rect 20700 4910 20920 4970
rect 20990 4910 21000 4970
rect 20700 4710 21000 4910
rect 20700 4650 20920 4710
rect 20990 4650 21000 4710
rect 20700 4450 21000 4650
rect 20700 4390 20920 4450
rect 20990 4390 21000 4450
rect 20700 4200 21000 4390
rect 21040 5350 21340 6300
rect 21040 5290 21050 5350
rect 21120 5290 21340 5350
rect 21040 5100 21340 5290
rect 21040 5030 21050 5100
rect 21120 5030 21340 5100
rect 21040 4840 21340 5030
rect 21040 4780 21050 4840
rect 21120 4780 21340 4840
rect 21040 4580 21340 4780
rect 21040 4520 21050 4580
rect 21120 4520 21340 4580
rect 21040 4320 21340 4520
rect 21040 4260 21050 4320
rect 21120 4260 21340 4320
rect 21040 4250 21130 4260
rect 20700 4160 20920 4200
rect 20370 4140 20920 4160
rect 20990 4140 21000 4200
rect 20290 3875 21000 4140
rect 20290 3865 20920 3875
rect 20290 3805 20300 3865
rect 20370 3855 20920 3865
rect 20370 3805 20590 3855
rect 20290 3615 20590 3805
rect 20290 3555 20300 3615
rect 20370 3555 20590 3615
rect 20290 3355 20590 3555
rect 20290 3295 20300 3355
rect 20370 3295 20590 3355
rect 20290 3105 20590 3295
rect 20290 3045 20300 3105
rect 20370 3045 20590 3105
rect 20290 2845 20590 3045
rect 20290 2785 20300 2845
rect 20370 2785 20590 2845
rect 20290 2585 20590 2785
rect 20290 2525 20300 2585
rect 20370 2525 20590 2585
rect 20290 2335 20590 2525
rect 20700 3815 20920 3855
rect 20990 3815 21000 3875
rect 20700 3625 21000 3815
rect 20700 3565 20920 3625
rect 20990 3565 21000 3625
rect 20700 3365 21000 3565
rect 20700 3305 20920 3365
rect 20990 3305 21000 3365
rect 20700 3105 21000 3305
rect 20700 3045 20920 3105
rect 20990 3045 21000 3105
rect 20700 2855 21000 3045
rect 20700 2795 20920 2855
rect 20990 2795 21000 2855
rect 20700 2595 21000 2795
rect 20700 2535 20920 2595
rect 20990 2535 21000 2595
rect 20700 2520 21000 2535
rect 21040 3755 21340 3765
rect 21040 3695 21050 3755
rect 21120 3695 21340 3755
rect 21040 3495 21340 3695
rect 21040 3435 21050 3495
rect 21120 3435 21340 3495
rect 21040 3235 21340 3435
rect 21040 3175 21050 3235
rect 21120 3175 21340 3235
rect 21040 2985 21340 3175
rect 21040 2915 21050 2985
rect 21120 2915 21340 2985
rect 21040 2725 21340 2915
rect 21040 2665 21050 2725
rect 21120 2665 21340 2725
rect 20290 2275 20300 2335
rect 20370 2275 20590 2335
rect 20290 2075 20590 2275
rect 20290 2015 20300 2075
rect 20370 2015 20590 2075
rect 20290 1855 20590 2015
rect 19200 1805 19770 1840
rect 18500 1620 18510 1690
rect 18570 1620 19100 1690
rect 18500 1430 19100 1620
rect 18500 1360 18510 1430
rect 18570 1360 19100 1430
rect 18500 1180 19100 1360
rect 21040 1310 21340 2665
rect 18500 1110 18510 1180
rect 18570 1110 19100 1180
rect 18500 920 19100 1110
rect 18500 850 18510 920
rect 18570 850 19100 920
rect 19240 1280 21340 1310
rect 19750 910 21340 1280
rect 19240 880 21340 910
rect 18500 670 19100 850
rect 18500 600 18510 670
rect 18570 600 19100 670
rect 17190 340 17720 410
rect 17780 340 17790 410
rect 17190 285 17790 340
rect 18500 410 19100 600
rect 18500 340 18510 410
rect 18570 340 19100 410
rect 18500 285 19100 340
rect 16970 -130 18090 285
rect 16970 -185 17400 -130
rect 17480 -135 17995 -130
rect 17480 -185 17785 -135
rect 16970 -190 17785 -185
rect 17865 -185 17995 -135
rect 18075 -185 18090 -130
rect 17865 -190 18090 -185
rect 16970 -250 18090 -190
rect 16970 -305 17080 -250
rect 17135 -305 17270 -250
rect 17325 -305 17465 -250
rect 17520 -305 17655 -250
rect 17710 -305 17850 -250
rect 17905 -305 18090 -250
rect 16970 -315 18090 -305
rect 18195 -40 20515 285
rect 18195 -240 19315 -40
rect 18195 -250 19320 -240
rect 18195 -305 18385 -250
rect 18440 -305 18580 -250
rect 18635 -305 18770 -250
rect 18825 -305 18965 -250
rect 19020 -305 19155 -250
rect 19210 -305 19320 -250
rect 18195 -315 19320 -305
rect 16965 -375 19765 -365
rect 16965 -430 16980 -375
rect 17035 -430 17175 -375
rect 17230 -430 17370 -375
rect 17425 -430 17560 -375
rect 17615 -430 17750 -375
rect 17805 -430 17945 -375
rect 18000 -430 18290 -375
rect 18345 -430 18485 -375
rect 18540 -430 18675 -375
rect 18730 -430 18865 -375
rect 18920 -430 19060 -375
rect 19115 -390 19255 -375
rect 19310 -390 19765 -375
rect 19115 -430 19230 -390
rect 16965 -940 19230 -430
rect 19730 -940 19765 -390
rect 16965 -965 19765 -940
<< via2 >>
rect 17450 7150 17705 7265
rect 18105 7150 18360 7265
rect 18750 7150 19005 7265
rect 19970 6120 20230 6135
rect 19970 6060 20170 6120
rect 20170 6060 20230 6120
rect 19970 5925 20230 6060
rect 19235 1840 19725 2215
rect 19230 -430 19255 -390
rect 19255 -430 19310 -390
rect 19310 -430 19730 -390
rect 19230 -940 19730 -430
<< metal3 >>
rect 17440 7265 20250 7275
rect 17440 7150 17450 7265
rect 17705 7150 18105 7265
rect 18360 7150 18750 7265
rect 19005 7150 20250 7265
rect 17440 7140 20250 7150
rect 19950 6135 20250 7140
rect 19950 5925 19970 6135
rect 20230 5925 20250 6135
rect 19950 5905 20250 5925
rect 19200 2215 19770 2255
rect 19200 1840 19235 2215
rect 19725 1840 19770 2215
rect 19200 1805 19770 1840
rect 19200 -390 19765 1805
rect 19200 -940 19230 -390
rect 19730 -940 19765 -390
rect 19200 -965 19765 -940
use sky130_fd_pr__pfet_01v8_lvt_D3M934  XM1
timestamp 1662404926
transform 0 1 20269 -1 0 2877
box -1127 -319 1127 319
use sky130_fd_pr__pfet_01v8_lvt_D3M934  XM2
timestamp 1662404926
transform 0 1 18069 -1 0 6117
box -1127 -319 1127 319
use sky130_fd_pr__pfet_01v8_lvt_D3M934  XM3
timestamp 1662404926
transform 0 1 18719 -1 0 6117
box -1127 -319 1127 319
use sky130_fd_pr__pfet_01v8_lvt_D3M934  XM29
timestamp 1662404926
transform 0 1 20269 -1 0 5127
box -1127 -319 1127 319
use sky130_fd_pr__pfet_01v8_lvt_D3ZSZ4  XM30
timestamp 1662404926
transform 0 1 21019 -1 0 3207
box -807 -319 807 319
use sky130_fd_pr__pfet_01v8_lvt_D3ZSZ4  XM31
timestamp 1662404926
transform 0 1 21019 -1 0 4807
box -807 -319 807 319
use sky130_fd_pr__pfet_01v8_lvt_D3M934  XM36
timestamp 1662404926
transform 0 1 17419 -1 0 6117
box -1127 -319 1127 319
use sky130_fd_pr__pfet_01v8_lvt_D3Z634  XM37
timestamp 1662404926
transform 0 1 17819 -1 0 2297
box -2087 -319 2087 319
use sky130_fd_pr__pfet_01v8_lvt_D3Z634  XM38
timestamp 1662404926
transform 0 1 18469 -1 0 2297
box -2087 -319 2087 319
use sky130_fd_pr__nfet_01v8_lvt_9DHFGX  XM39
timestamp 1662404926
transform 1 0 17493 0 1 -340
box -647 -310 647 310
use sky130_fd_pr__nfet_01v8_lvt_9DHFGX  XM40
timestamp 1662404926
transform -1 0 18797 0 -1 -340
box -647 -310 647 310
use sky130_fd_pr__res_high_po_2p85_P79JE3  XR19
timestamp 1662404926
transform 1 0 19491 0 1 5548
box -451 -1358 451 1358
use sky130_fd_pr__res_high_po_2p85_MM89SS  XR20
timestamp 1662404926
transform 1 0 19491 0 1 2448
box -451 -1738 451 1738
<< labels >>
rlabel metal1 20820 5520 21340 5580 1 AMP
rlabel metal1 21020 2435 21340 2495 1 VOP
rlabel metal3 18360 7140 18750 7275 1 VDD
rlabel metal2 19060 -40 20515 285 1 BIASOUT
rlabel locali 18970 6975 20025 7020 1 PSUB
rlabel metal1 17220 7150 20470 7220 1 BIAS2V
rlabel metal1 17100 4310 18020 4370 1 VCTRL
rlabel metal2 16965 -965 19230 -430 1 GND
rlabel locali 19070 -100 19115 790 1 SUB
<< end >>
