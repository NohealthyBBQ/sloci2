magic
tech sky130A
timestamp 1671727289
<< metal1 >>
rect 525 790 530 850
rect 560 790 565 850
rect 0 350 130 360
rect -95 320 -90 350
rect -60 320 -55 350
rect 0 320 10 350
rect 40 320 130 350
rect 675 320 680 350
rect 710 320 715 350
rect 0 310 130 320
rect 295 250 300 280
rect 330 250 335 280
rect 865 250 870 280
rect 900 250 905 280
rect 525 -170 530 -110
rect 560 -170 565 -110
rect 105 -560 110 -530
rect 140 -560 145 -530
rect 675 -560 680 -530
rect 710 -560 715 -530
rect 5 -640 10 -610
rect 40 -640 45 -610
rect -85 -720 -80 -690
rect -50 -720 -45 -690
rect 295 -720 300 -690
rect 330 -720 335 -690
rect 865 -720 870 -690
rect 900 -720 905 -690
<< via1 >>
rect 530 790 560 850
rect -90 320 -60 350
rect 10 320 40 350
rect 680 320 710 350
rect 300 250 330 280
rect 870 250 900 280
rect 530 -170 560 -110
rect 110 -560 140 -530
rect 680 -560 710 -530
rect 10 -640 40 -610
rect -80 -720 -50 -690
rect 300 -720 330 -690
rect 870 -720 900 -690
<< metal2 >>
rect 530 850 1180 860
rect 560 790 1180 850
rect 530 780 1180 790
rect -90 520 710 550
rect -90 350 -60 520
rect -90 40 -60 320
rect 10 350 40 360
rect 10 40 40 320
rect 680 350 710 520
rect 680 310 710 320
rect 300 280 330 285
rect 870 280 900 285
rect 330 250 440 280
rect 300 245 330 250
rect 300 40 330 45
rect 10 10 140 40
rect -90 0 -60 10
rect 10 -40 40 -35
rect 10 -610 40 -70
rect 110 -530 140 10
rect 300 -530 330 10
rect 410 -40 440 250
rect 900 250 1010 280
rect 870 245 900 250
rect 410 -80 440 -70
rect 980 -40 1010 250
rect 980 -75 1010 -70
rect 530 -110 1180 -100
rect 560 -170 1180 -110
rect 530 -180 1180 -170
rect 680 -530 710 -525
rect 300 -560 680 -530
rect 110 -565 140 -560
rect 680 -565 710 -560
rect 10 -650 40 -640
rect -80 -690 -50 -685
rect 300 -690 330 -685
rect 870 -690 900 -685
rect -50 -720 300 -690
rect 330 -720 870 -690
rect -80 -725 -50 -720
rect 300 -725 330 -720
rect 870 -725 900 -720
<< via2 >>
rect -90 10 -60 40
rect 10 -70 40 -40
rect 300 10 330 40
rect 410 -70 440 -40
rect 980 -70 1010 -40
<< metal3 >>
rect -110 40 340 50
rect -110 10 -90 40
rect -60 10 300 40
rect 330 10 340 40
rect -110 0 340 10
rect 0 -40 1030 -30
rect 0 -70 10 -40
rect 40 -70 410 -40
rect 440 -70 980 -40
rect 1010 -70 1030 -40
rect 0 -80 1030 -70
use and  and_0
timestamp 1671683902
transform 1 0 580 0 1 -630
box -10 -330 616 594
use and  and_1
timestamp 1671683902
transform 1 0 10 0 1 -630
box -10 -330 616 594
use and  and_2
timestamp 1671683902
transform 1 0 580 0 1 330
box -10 -330 616 594
use and  and_3
timestamp 1671683902
transform 1 0 10 0 1 330
box -10 -330 616 594
use inv  inv_0
timestamp 1671682090
transform 1 0 -160 0 1 -580
box -30 -380 216 544
use inv  inv_1
timestamp 1671682090
transform 1 0 -160 0 1 380
box -30 -380 216 544
<< labels >>
flabel space 0 310 135 360 0 FreeSans 320 0 0 0 A_b
flabel metal2 10 -610 40 -70 0 FreeSans 320 0 0 0 B_b
<< end >>
