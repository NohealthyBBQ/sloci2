magic
tech sky130A
magscale 1 2
timestamp 1671675948
<< nwell >>
rect -246 -419 246 419
<< pmos >>
rect -50 -200 50 200
<< pdiff >>
rect -108 188 -50 200
rect -108 -188 -96 188
rect -62 -188 -50 188
rect -108 -200 -50 -188
rect 50 188 108 200
rect 50 -188 62 188
rect 96 -188 108 188
rect 50 -200 108 -188
<< pdiffc >>
rect -96 -188 -62 188
rect 62 -188 96 188
<< nsubdiff >>
rect -210 349 -114 383
rect 114 349 210 383
rect -210 287 -176 349
rect 176 287 210 349
rect -210 -349 -176 -287
rect 176 -349 210 -287
rect -210 -383 -114 -349
rect 114 -383 210 -349
<< nsubdiffcont >>
rect -114 349 114 383
rect -210 -287 -176 287
rect 176 -287 210 287
rect -114 -383 114 -349
<< poly >>
rect -50 281 50 297
rect -50 247 -34 281
rect 34 247 50 281
rect -50 200 50 247
rect -50 -247 50 -200
rect -50 -281 -34 -247
rect 34 -281 50 -247
rect -50 -297 50 -281
<< polycont >>
rect -34 247 34 281
rect -34 -281 34 -247
<< locali >>
rect -210 349 -114 383
rect 114 349 210 383
rect -210 287 -176 349
rect 176 287 210 349
rect -50 247 -34 281
rect 34 247 50 281
rect -96 188 -62 204
rect -96 -204 -62 -188
rect 62 188 96 204
rect 62 -204 96 -188
rect -50 -281 -34 -247
rect 34 -281 50 -247
rect -210 -349 -176 -287
rect 176 -349 210 -287
rect -210 -383 -114 -349
rect 114 -383 210 -349
<< viali >>
rect -34 247 34 281
rect -96 -188 -62 188
rect 62 -188 96 188
rect -34 -281 34 -247
<< metal1 >>
rect -46 281 46 287
rect -46 247 -34 281
rect 34 247 46 281
rect -46 241 46 247
rect -102 188 -56 200
rect -102 -188 -96 188
rect -62 -188 -56 188
rect -102 -200 -56 -188
rect 56 188 102 200
rect 56 -188 62 188
rect 96 -188 102 188
rect 56 -200 102 -188
rect -46 -247 46 -241
rect -46 -281 -34 -247
rect 34 -281 46 -247
rect -46 -287 46 -281
<< properties >>
string FIXED_BBOX -193 -366 193 366
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 2 l 0.5 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
