magic
tech sky130A
magscale 1 2
timestamp 1662732419
<< metal3 >>
rect -1750 -2100 1620 2100
<< mimcap >>
rect -1650 1960 1550 2000
rect -1650 -1960 -1610 1960
rect 1510 -1960 1550 1960
rect -1650 -2000 1550 -1960
<< mimcapcontact >>
rect -1610 -1960 1510 1960
<< metal4 >>
rect -1611 1960 1511 1961
rect -1611 -1960 -1610 1960
rect 1510 -1960 1511 1960
rect -1611 -1961 1511 -1960
<< properties >>
string FIXED_BBOX -1750 -2100 1650 2100
string gencell sky130_fd_pr__cap_mim_m3_1
string library sky130
string parameters w 16 l 20 val 653.68 carea 2.00 cperi 0.19 nx 1 ny 1 dummy 0 square 0 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 1 tconnect 1 ccov 100
<< end >>
