magic
tech sky130A
magscale 1 2
timestamp 1662407989
<< error_p >>
rect -2765 172 -2707 178
rect -2573 172 -2515 178
rect -2381 172 -2323 178
rect -2189 172 -2131 178
rect -1997 172 -1939 178
rect -1805 172 -1747 178
rect -1613 172 -1555 178
rect -1421 172 -1363 178
rect -1229 172 -1171 178
rect -1037 172 -979 178
rect -845 172 -787 178
rect -653 172 -595 178
rect -461 172 -403 178
rect -269 172 -211 178
rect -77 172 -19 178
rect 115 172 173 178
rect 307 172 365 178
rect 499 172 557 178
rect 691 172 749 178
rect 883 172 941 178
rect 1075 172 1133 178
rect 1267 172 1325 178
rect 1459 172 1517 178
rect 1651 172 1709 178
rect 1843 172 1901 178
rect 2035 172 2093 178
rect 2227 172 2285 178
rect 2419 172 2477 178
rect 2611 172 2669 178
rect 2803 172 2861 178
rect -2765 138 -2753 172
rect -2573 138 -2561 172
rect -2381 138 -2369 172
rect -2189 138 -2177 172
rect -1997 138 -1985 172
rect -1805 138 -1793 172
rect -1613 138 -1601 172
rect -1421 138 -1409 172
rect -1229 138 -1217 172
rect -1037 138 -1025 172
rect -845 138 -833 172
rect -653 138 -641 172
rect -461 138 -449 172
rect -269 138 -257 172
rect -77 138 -65 172
rect 115 138 127 172
rect 307 138 319 172
rect 499 138 511 172
rect 691 138 703 172
rect 883 138 895 172
rect 1075 138 1087 172
rect 1267 138 1279 172
rect 1459 138 1471 172
rect 1651 138 1663 172
rect 1843 138 1855 172
rect 2035 138 2047 172
rect 2227 138 2239 172
rect 2419 138 2431 172
rect 2611 138 2623 172
rect 2803 138 2815 172
rect -2765 132 -2707 138
rect -2573 132 -2515 138
rect -2381 132 -2323 138
rect -2189 132 -2131 138
rect -1997 132 -1939 138
rect -1805 132 -1747 138
rect -1613 132 -1555 138
rect -1421 132 -1363 138
rect -1229 132 -1171 138
rect -1037 132 -979 138
rect -845 132 -787 138
rect -653 132 -595 138
rect -461 132 -403 138
rect -269 132 -211 138
rect -77 132 -19 138
rect 115 132 173 138
rect 307 132 365 138
rect 499 132 557 138
rect 691 132 749 138
rect 883 132 941 138
rect 1075 132 1133 138
rect 1267 132 1325 138
rect 1459 132 1517 138
rect 1651 132 1709 138
rect 1843 132 1901 138
rect 2035 132 2093 138
rect 2227 132 2285 138
rect 2419 132 2477 138
rect 2611 132 2669 138
rect 2803 132 2861 138
rect -2861 -138 -2803 -132
rect -2669 -138 -2611 -132
rect -2477 -138 -2419 -132
rect -2285 -138 -2227 -132
rect -2093 -138 -2035 -132
rect -1901 -138 -1843 -132
rect -1709 -138 -1651 -132
rect -1517 -138 -1459 -132
rect -1325 -138 -1267 -132
rect -1133 -138 -1075 -132
rect -941 -138 -883 -132
rect -749 -138 -691 -132
rect -557 -138 -499 -132
rect -365 -138 -307 -132
rect -173 -138 -115 -132
rect 19 -138 77 -132
rect 211 -138 269 -132
rect 403 -138 461 -132
rect 595 -138 653 -132
rect 787 -138 845 -132
rect 979 -138 1037 -132
rect 1171 -138 1229 -132
rect 1363 -138 1421 -132
rect 1555 -138 1613 -132
rect 1747 -138 1805 -132
rect 1939 -138 1997 -132
rect 2131 -138 2189 -132
rect 2323 -138 2381 -132
rect 2515 -138 2573 -132
rect 2707 -138 2765 -132
rect -2861 -172 -2849 -138
rect -2669 -172 -2657 -138
rect -2477 -172 -2465 -138
rect -2285 -172 -2273 -138
rect -2093 -172 -2081 -138
rect -1901 -172 -1889 -138
rect -1709 -172 -1697 -138
rect -1517 -172 -1505 -138
rect -1325 -172 -1313 -138
rect -1133 -172 -1121 -138
rect -941 -172 -929 -138
rect -749 -172 -737 -138
rect -557 -172 -545 -138
rect -365 -172 -353 -138
rect -173 -172 -161 -138
rect 19 -172 31 -138
rect 211 -172 223 -138
rect 403 -172 415 -138
rect 595 -172 607 -138
rect 787 -172 799 -138
rect 979 -172 991 -138
rect 1171 -172 1183 -138
rect 1363 -172 1375 -138
rect 1555 -172 1567 -138
rect 1747 -172 1759 -138
rect 1939 -172 1951 -138
rect 2131 -172 2143 -138
rect 2323 -172 2335 -138
rect 2515 -172 2527 -138
rect 2707 -172 2719 -138
rect -2861 -178 -2803 -172
rect -2669 -178 -2611 -172
rect -2477 -178 -2419 -172
rect -2285 -178 -2227 -172
rect -2093 -178 -2035 -172
rect -1901 -178 -1843 -172
rect -1709 -178 -1651 -172
rect -1517 -178 -1459 -172
rect -1325 -178 -1267 -172
rect -1133 -178 -1075 -172
rect -941 -178 -883 -172
rect -749 -178 -691 -172
rect -557 -178 -499 -172
rect -365 -178 -307 -172
rect -173 -178 -115 -172
rect 19 -178 77 -172
rect 211 -178 269 -172
rect 403 -178 461 -172
rect 595 -178 653 -172
rect 787 -178 845 -172
rect 979 -178 1037 -172
rect 1171 -178 1229 -172
rect 1363 -178 1421 -172
rect 1555 -178 1613 -172
rect 1747 -178 1805 -172
rect 1939 -178 1997 -172
rect 2131 -178 2189 -172
rect 2323 -178 2381 -172
rect 2515 -178 2573 -172
rect 2707 -178 2765 -172
<< pwell >>
rect -3047 -310 3047 310
<< nmoslvt >>
rect -2847 -100 -2817 100
rect -2751 -100 -2721 100
rect -2655 -100 -2625 100
rect -2559 -100 -2529 100
rect -2463 -100 -2433 100
rect -2367 -100 -2337 100
rect -2271 -100 -2241 100
rect -2175 -100 -2145 100
rect -2079 -100 -2049 100
rect -1983 -100 -1953 100
rect -1887 -100 -1857 100
rect -1791 -100 -1761 100
rect -1695 -100 -1665 100
rect -1599 -100 -1569 100
rect -1503 -100 -1473 100
rect -1407 -100 -1377 100
rect -1311 -100 -1281 100
rect -1215 -100 -1185 100
rect -1119 -100 -1089 100
rect -1023 -100 -993 100
rect -927 -100 -897 100
rect -831 -100 -801 100
rect -735 -100 -705 100
rect -639 -100 -609 100
rect -543 -100 -513 100
rect -447 -100 -417 100
rect -351 -100 -321 100
rect -255 -100 -225 100
rect -159 -100 -129 100
rect -63 -100 -33 100
rect 33 -100 63 100
rect 129 -100 159 100
rect 225 -100 255 100
rect 321 -100 351 100
rect 417 -100 447 100
rect 513 -100 543 100
rect 609 -100 639 100
rect 705 -100 735 100
rect 801 -100 831 100
rect 897 -100 927 100
rect 993 -100 1023 100
rect 1089 -100 1119 100
rect 1185 -100 1215 100
rect 1281 -100 1311 100
rect 1377 -100 1407 100
rect 1473 -100 1503 100
rect 1569 -100 1599 100
rect 1665 -100 1695 100
rect 1761 -100 1791 100
rect 1857 -100 1887 100
rect 1953 -100 1983 100
rect 2049 -100 2079 100
rect 2145 -100 2175 100
rect 2241 -100 2271 100
rect 2337 -100 2367 100
rect 2433 -100 2463 100
rect 2529 -100 2559 100
rect 2625 -100 2655 100
rect 2721 -100 2751 100
rect 2817 -100 2847 100
<< ndiff >>
rect -2909 88 -2847 100
rect -2909 -88 -2897 88
rect -2863 -88 -2847 88
rect -2909 -100 -2847 -88
rect -2817 88 -2751 100
rect -2817 -88 -2801 88
rect -2767 -88 -2751 88
rect -2817 -100 -2751 -88
rect -2721 88 -2655 100
rect -2721 -88 -2705 88
rect -2671 -88 -2655 88
rect -2721 -100 -2655 -88
rect -2625 88 -2559 100
rect -2625 -88 -2609 88
rect -2575 -88 -2559 88
rect -2625 -100 -2559 -88
rect -2529 88 -2463 100
rect -2529 -88 -2513 88
rect -2479 -88 -2463 88
rect -2529 -100 -2463 -88
rect -2433 88 -2367 100
rect -2433 -88 -2417 88
rect -2383 -88 -2367 88
rect -2433 -100 -2367 -88
rect -2337 88 -2271 100
rect -2337 -88 -2321 88
rect -2287 -88 -2271 88
rect -2337 -100 -2271 -88
rect -2241 88 -2175 100
rect -2241 -88 -2225 88
rect -2191 -88 -2175 88
rect -2241 -100 -2175 -88
rect -2145 88 -2079 100
rect -2145 -88 -2129 88
rect -2095 -88 -2079 88
rect -2145 -100 -2079 -88
rect -2049 88 -1983 100
rect -2049 -88 -2033 88
rect -1999 -88 -1983 88
rect -2049 -100 -1983 -88
rect -1953 88 -1887 100
rect -1953 -88 -1937 88
rect -1903 -88 -1887 88
rect -1953 -100 -1887 -88
rect -1857 88 -1791 100
rect -1857 -88 -1841 88
rect -1807 -88 -1791 88
rect -1857 -100 -1791 -88
rect -1761 88 -1695 100
rect -1761 -88 -1745 88
rect -1711 -88 -1695 88
rect -1761 -100 -1695 -88
rect -1665 88 -1599 100
rect -1665 -88 -1649 88
rect -1615 -88 -1599 88
rect -1665 -100 -1599 -88
rect -1569 88 -1503 100
rect -1569 -88 -1553 88
rect -1519 -88 -1503 88
rect -1569 -100 -1503 -88
rect -1473 88 -1407 100
rect -1473 -88 -1457 88
rect -1423 -88 -1407 88
rect -1473 -100 -1407 -88
rect -1377 88 -1311 100
rect -1377 -88 -1361 88
rect -1327 -88 -1311 88
rect -1377 -100 -1311 -88
rect -1281 88 -1215 100
rect -1281 -88 -1265 88
rect -1231 -88 -1215 88
rect -1281 -100 -1215 -88
rect -1185 88 -1119 100
rect -1185 -88 -1169 88
rect -1135 -88 -1119 88
rect -1185 -100 -1119 -88
rect -1089 88 -1023 100
rect -1089 -88 -1073 88
rect -1039 -88 -1023 88
rect -1089 -100 -1023 -88
rect -993 88 -927 100
rect -993 -88 -977 88
rect -943 -88 -927 88
rect -993 -100 -927 -88
rect -897 88 -831 100
rect -897 -88 -881 88
rect -847 -88 -831 88
rect -897 -100 -831 -88
rect -801 88 -735 100
rect -801 -88 -785 88
rect -751 -88 -735 88
rect -801 -100 -735 -88
rect -705 88 -639 100
rect -705 -88 -689 88
rect -655 -88 -639 88
rect -705 -100 -639 -88
rect -609 88 -543 100
rect -609 -88 -593 88
rect -559 -88 -543 88
rect -609 -100 -543 -88
rect -513 88 -447 100
rect -513 -88 -497 88
rect -463 -88 -447 88
rect -513 -100 -447 -88
rect -417 88 -351 100
rect -417 -88 -401 88
rect -367 -88 -351 88
rect -417 -100 -351 -88
rect -321 88 -255 100
rect -321 -88 -305 88
rect -271 -88 -255 88
rect -321 -100 -255 -88
rect -225 88 -159 100
rect -225 -88 -209 88
rect -175 -88 -159 88
rect -225 -100 -159 -88
rect -129 88 -63 100
rect -129 -88 -113 88
rect -79 -88 -63 88
rect -129 -100 -63 -88
rect -33 88 33 100
rect -33 -88 -17 88
rect 17 -88 33 88
rect -33 -100 33 -88
rect 63 88 129 100
rect 63 -88 79 88
rect 113 -88 129 88
rect 63 -100 129 -88
rect 159 88 225 100
rect 159 -88 175 88
rect 209 -88 225 88
rect 159 -100 225 -88
rect 255 88 321 100
rect 255 -88 271 88
rect 305 -88 321 88
rect 255 -100 321 -88
rect 351 88 417 100
rect 351 -88 367 88
rect 401 -88 417 88
rect 351 -100 417 -88
rect 447 88 513 100
rect 447 -88 463 88
rect 497 -88 513 88
rect 447 -100 513 -88
rect 543 88 609 100
rect 543 -88 559 88
rect 593 -88 609 88
rect 543 -100 609 -88
rect 639 88 705 100
rect 639 -88 655 88
rect 689 -88 705 88
rect 639 -100 705 -88
rect 735 88 801 100
rect 735 -88 751 88
rect 785 -88 801 88
rect 735 -100 801 -88
rect 831 88 897 100
rect 831 -88 847 88
rect 881 -88 897 88
rect 831 -100 897 -88
rect 927 88 993 100
rect 927 -88 943 88
rect 977 -88 993 88
rect 927 -100 993 -88
rect 1023 88 1089 100
rect 1023 -88 1039 88
rect 1073 -88 1089 88
rect 1023 -100 1089 -88
rect 1119 88 1185 100
rect 1119 -88 1135 88
rect 1169 -88 1185 88
rect 1119 -100 1185 -88
rect 1215 88 1281 100
rect 1215 -88 1231 88
rect 1265 -88 1281 88
rect 1215 -100 1281 -88
rect 1311 88 1377 100
rect 1311 -88 1327 88
rect 1361 -88 1377 88
rect 1311 -100 1377 -88
rect 1407 88 1473 100
rect 1407 -88 1423 88
rect 1457 -88 1473 88
rect 1407 -100 1473 -88
rect 1503 88 1569 100
rect 1503 -88 1519 88
rect 1553 -88 1569 88
rect 1503 -100 1569 -88
rect 1599 88 1665 100
rect 1599 -88 1615 88
rect 1649 -88 1665 88
rect 1599 -100 1665 -88
rect 1695 88 1761 100
rect 1695 -88 1711 88
rect 1745 -88 1761 88
rect 1695 -100 1761 -88
rect 1791 88 1857 100
rect 1791 -88 1807 88
rect 1841 -88 1857 88
rect 1791 -100 1857 -88
rect 1887 88 1953 100
rect 1887 -88 1903 88
rect 1937 -88 1953 88
rect 1887 -100 1953 -88
rect 1983 88 2049 100
rect 1983 -88 1999 88
rect 2033 -88 2049 88
rect 1983 -100 2049 -88
rect 2079 88 2145 100
rect 2079 -88 2095 88
rect 2129 -88 2145 88
rect 2079 -100 2145 -88
rect 2175 88 2241 100
rect 2175 -88 2191 88
rect 2225 -88 2241 88
rect 2175 -100 2241 -88
rect 2271 88 2337 100
rect 2271 -88 2287 88
rect 2321 -88 2337 88
rect 2271 -100 2337 -88
rect 2367 88 2433 100
rect 2367 -88 2383 88
rect 2417 -88 2433 88
rect 2367 -100 2433 -88
rect 2463 88 2529 100
rect 2463 -88 2479 88
rect 2513 -88 2529 88
rect 2463 -100 2529 -88
rect 2559 88 2625 100
rect 2559 -88 2575 88
rect 2609 -88 2625 88
rect 2559 -100 2625 -88
rect 2655 88 2721 100
rect 2655 -88 2671 88
rect 2705 -88 2721 88
rect 2655 -100 2721 -88
rect 2751 88 2817 100
rect 2751 -88 2767 88
rect 2801 -88 2817 88
rect 2751 -100 2817 -88
rect 2847 88 2909 100
rect 2847 -88 2863 88
rect 2897 -88 2909 88
rect 2847 -100 2909 -88
<< ndiffc >>
rect -2897 -88 -2863 88
rect -2801 -88 -2767 88
rect -2705 -88 -2671 88
rect -2609 -88 -2575 88
rect -2513 -88 -2479 88
rect -2417 -88 -2383 88
rect -2321 -88 -2287 88
rect -2225 -88 -2191 88
rect -2129 -88 -2095 88
rect -2033 -88 -1999 88
rect -1937 -88 -1903 88
rect -1841 -88 -1807 88
rect -1745 -88 -1711 88
rect -1649 -88 -1615 88
rect -1553 -88 -1519 88
rect -1457 -88 -1423 88
rect -1361 -88 -1327 88
rect -1265 -88 -1231 88
rect -1169 -88 -1135 88
rect -1073 -88 -1039 88
rect -977 -88 -943 88
rect -881 -88 -847 88
rect -785 -88 -751 88
rect -689 -88 -655 88
rect -593 -88 -559 88
rect -497 -88 -463 88
rect -401 -88 -367 88
rect -305 -88 -271 88
rect -209 -88 -175 88
rect -113 -88 -79 88
rect -17 -88 17 88
rect 79 -88 113 88
rect 175 -88 209 88
rect 271 -88 305 88
rect 367 -88 401 88
rect 463 -88 497 88
rect 559 -88 593 88
rect 655 -88 689 88
rect 751 -88 785 88
rect 847 -88 881 88
rect 943 -88 977 88
rect 1039 -88 1073 88
rect 1135 -88 1169 88
rect 1231 -88 1265 88
rect 1327 -88 1361 88
rect 1423 -88 1457 88
rect 1519 -88 1553 88
rect 1615 -88 1649 88
rect 1711 -88 1745 88
rect 1807 -88 1841 88
rect 1903 -88 1937 88
rect 1999 -88 2033 88
rect 2095 -88 2129 88
rect 2191 -88 2225 88
rect 2287 -88 2321 88
rect 2383 -88 2417 88
rect 2479 -88 2513 88
rect 2575 -88 2609 88
rect 2671 -88 2705 88
rect 2767 -88 2801 88
rect 2863 -88 2897 88
<< psubdiff >>
rect -3011 240 -2915 274
rect 2915 240 3011 274
rect -3011 178 -2977 240
rect 2977 178 3011 240
rect -3011 -240 -2977 -178
rect 2977 -240 3011 -178
rect -3011 -274 -2915 -240
rect 2915 -274 3011 -240
<< psubdiffcont >>
rect -2915 240 2915 274
rect -3011 -178 -2977 178
rect 2977 -178 3011 178
rect -2915 -274 2915 -240
<< poly >>
rect -2769 172 -2703 188
rect -2769 138 -2753 172
rect -2719 138 -2703 172
rect -2847 100 -2817 126
rect -2769 122 -2703 138
rect -2577 172 -2511 188
rect -2577 138 -2561 172
rect -2527 138 -2511 172
rect -2751 100 -2721 122
rect -2655 100 -2625 126
rect -2577 122 -2511 138
rect -2385 172 -2319 188
rect -2385 138 -2369 172
rect -2335 138 -2319 172
rect -2559 100 -2529 122
rect -2463 100 -2433 126
rect -2385 122 -2319 138
rect -2193 172 -2127 188
rect -2193 138 -2177 172
rect -2143 138 -2127 172
rect -2367 100 -2337 122
rect -2271 100 -2241 126
rect -2193 122 -2127 138
rect -2001 172 -1935 188
rect -2001 138 -1985 172
rect -1951 138 -1935 172
rect -2175 100 -2145 122
rect -2079 100 -2049 126
rect -2001 122 -1935 138
rect -1809 172 -1743 188
rect -1809 138 -1793 172
rect -1759 138 -1743 172
rect -1983 100 -1953 122
rect -1887 100 -1857 126
rect -1809 122 -1743 138
rect -1617 172 -1551 188
rect -1617 138 -1601 172
rect -1567 138 -1551 172
rect -1791 100 -1761 122
rect -1695 100 -1665 126
rect -1617 122 -1551 138
rect -1425 172 -1359 188
rect -1425 138 -1409 172
rect -1375 138 -1359 172
rect -1599 100 -1569 122
rect -1503 100 -1473 126
rect -1425 122 -1359 138
rect -1233 172 -1167 188
rect -1233 138 -1217 172
rect -1183 138 -1167 172
rect -1407 100 -1377 122
rect -1311 100 -1281 126
rect -1233 122 -1167 138
rect -1041 172 -975 188
rect -1041 138 -1025 172
rect -991 138 -975 172
rect -1215 100 -1185 122
rect -1119 100 -1089 126
rect -1041 122 -975 138
rect -849 172 -783 188
rect -849 138 -833 172
rect -799 138 -783 172
rect -1023 100 -993 122
rect -927 100 -897 126
rect -849 122 -783 138
rect -657 172 -591 188
rect -657 138 -641 172
rect -607 138 -591 172
rect -831 100 -801 122
rect -735 100 -705 126
rect -657 122 -591 138
rect -465 172 -399 188
rect -465 138 -449 172
rect -415 138 -399 172
rect -639 100 -609 122
rect -543 100 -513 126
rect -465 122 -399 138
rect -273 172 -207 188
rect -273 138 -257 172
rect -223 138 -207 172
rect -447 100 -417 122
rect -351 100 -321 126
rect -273 122 -207 138
rect -81 172 -15 188
rect -81 138 -65 172
rect -31 138 -15 172
rect -255 100 -225 122
rect -159 100 -129 126
rect -81 122 -15 138
rect 111 172 177 188
rect 111 138 127 172
rect 161 138 177 172
rect -63 100 -33 122
rect 33 100 63 126
rect 111 122 177 138
rect 303 172 369 188
rect 303 138 319 172
rect 353 138 369 172
rect 129 100 159 122
rect 225 100 255 126
rect 303 122 369 138
rect 495 172 561 188
rect 495 138 511 172
rect 545 138 561 172
rect 321 100 351 122
rect 417 100 447 126
rect 495 122 561 138
rect 687 172 753 188
rect 687 138 703 172
rect 737 138 753 172
rect 513 100 543 122
rect 609 100 639 126
rect 687 122 753 138
rect 879 172 945 188
rect 879 138 895 172
rect 929 138 945 172
rect 705 100 735 122
rect 801 100 831 126
rect 879 122 945 138
rect 1071 172 1137 188
rect 1071 138 1087 172
rect 1121 138 1137 172
rect 897 100 927 122
rect 993 100 1023 126
rect 1071 122 1137 138
rect 1263 172 1329 188
rect 1263 138 1279 172
rect 1313 138 1329 172
rect 1089 100 1119 122
rect 1185 100 1215 126
rect 1263 122 1329 138
rect 1455 172 1521 188
rect 1455 138 1471 172
rect 1505 138 1521 172
rect 1281 100 1311 122
rect 1377 100 1407 126
rect 1455 122 1521 138
rect 1647 172 1713 188
rect 1647 138 1663 172
rect 1697 138 1713 172
rect 1473 100 1503 122
rect 1569 100 1599 126
rect 1647 122 1713 138
rect 1839 172 1905 188
rect 1839 138 1855 172
rect 1889 138 1905 172
rect 1665 100 1695 122
rect 1761 100 1791 126
rect 1839 122 1905 138
rect 2031 172 2097 188
rect 2031 138 2047 172
rect 2081 138 2097 172
rect 1857 100 1887 122
rect 1953 100 1983 126
rect 2031 122 2097 138
rect 2223 172 2289 188
rect 2223 138 2239 172
rect 2273 138 2289 172
rect 2049 100 2079 122
rect 2145 100 2175 126
rect 2223 122 2289 138
rect 2415 172 2481 188
rect 2415 138 2431 172
rect 2465 138 2481 172
rect 2241 100 2271 122
rect 2337 100 2367 126
rect 2415 122 2481 138
rect 2607 172 2673 188
rect 2607 138 2623 172
rect 2657 138 2673 172
rect 2433 100 2463 122
rect 2529 100 2559 126
rect 2607 122 2673 138
rect 2799 172 2865 188
rect 2799 138 2815 172
rect 2849 138 2865 172
rect 2625 100 2655 122
rect 2721 100 2751 126
rect 2799 122 2865 138
rect 2817 100 2847 122
rect -2847 -122 -2817 -100
rect -2865 -138 -2799 -122
rect -2751 -126 -2721 -100
rect -2655 -122 -2625 -100
rect -2865 -172 -2849 -138
rect -2815 -172 -2799 -138
rect -2865 -188 -2799 -172
rect -2673 -138 -2607 -122
rect -2559 -126 -2529 -100
rect -2463 -122 -2433 -100
rect -2673 -172 -2657 -138
rect -2623 -172 -2607 -138
rect -2673 -188 -2607 -172
rect -2481 -138 -2415 -122
rect -2367 -126 -2337 -100
rect -2271 -122 -2241 -100
rect -2481 -172 -2465 -138
rect -2431 -172 -2415 -138
rect -2481 -188 -2415 -172
rect -2289 -138 -2223 -122
rect -2175 -126 -2145 -100
rect -2079 -122 -2049 -100
rect -2289 -172 -2273 -138
rect -2239 -172 -2223 -138
rect -2289 -188 -2223 -172
rect -2097 -138 -2031 -122
rect -1983 -126 -1953 -100
rect -1887 -122 -1857 -100
rect -2097 -172 -2081 -138
rect -2047 -172 -2031 -138
rect -2097 -188 -2031 -172
rect -1905 -138 -1839 -122
rect -1791 -126 -1761 -100
rect -1695 -122 -1665 -100
rect -1905 -172 -1889 -138
rect -1855 -172 -1839 -138
rect -1905 -188 -1839 -172
rect -1713 -138 -1647 -122
rect -1599 -126 -1569 -100
rect -1503 -122 -1473 -100
rect -1713 -172 -1697 -138
rect -1663 -172 -1647 -138
rect -1713 -188 -1647 -172
rect -1521 -138 -1455 -122
rect -1407 -126 -1377 -100
rect -1311 -122 -1281 -100
rect -1521 -172 -1505 -138
rect -1471 -172 -1455 -138
rect -1521 -188 -1455 -172
rect -1329 -138 -1263 -122
rect -1215 -126 -1185 -100
rect -1119 -122 -1089 -100
rect -1329 -172 -1313 -138
rect -1279 -172 -1263 -138
rect -1329 -188 -1263 -172
rect -1137 -138 -1071 -122
rect -1023 -126 -993 -100
rect -927 -122 -897 -100
rect -1137 -172 -1121 -138
rect -1087 -172 -1071 -138
rect -1137 -188 -1071 -172
rect -945 -138 -879 -122
rect -831 -126 -801 -100
rect -735 -122 -705 -100
rect -945 -172 -929 -138
rect -895 -172 -879 -138
rect -945 -188 -879 -172
rect -753 -138 -687 -122
rect -639 -126 -609 -100
rect -543 -122 -513 -100
rect -753 -172 -737 -138
rect -703 -172 -687 -138
rect -753 -188 -687 -172
rect -561 -138 -495 -122
rect -447 -126 -417 -100
rect -351 -122 -321 -100
rect -561 -172 -545 -138
rect -511 -172 -495 -138
rect -561 -188 -495 -172
rect -369 -138 -303 -122
rect -255 -126 -225 -100
rect -159 -122 -129 -100
rect -369 -172 -353 -138
rect -319 -172 -303 -138
rect -369 -188 -303 -172
rect -177 -138 -111 -122
rect -63 -126 -33 -100
rect 33 -122 63 -100
rect -177 -172 -161 -138
rect -127 -172 -111 -138
rect -177 -188 -111 -172
rect 15 -138 81 -122
rect 129 -126 159 -100
rect 225 -122 255 -100
rect 15 -172 31 -138
rect 65 -172 81 -138
rect 15 -188 81 -172
rect 207 -138 273 -122
rect 321 -126 351 -100
rect 417 -122 447 -100
rect 207 -172 223 -138
rect 257 -172 273 -138
rect 207 -188 273 -172
rect 399 -138 465 -122
rect 513 -126 543 -100
rect 609 -122 639 -100
rect 399 -172 415 -138
rect 449 -172 465 -138
rect 399 -188 465 -172
rect 591 -138 657 -122
rect 705 -126 735 -100
rect 801 -122 831 -100
rect 591 -172 607 -138
rect 641 -172 657 -138
rect 591 -188 657 -172
rect 783 -138 849 -122
rect 897 -126 927 -100
rect 993 -122 1023 -100
rect 783 -172 799 -138
rect 833 -172 849 -138
rect 783 -188 849 -172
rect 975 -138 1041 -122
rect 1089 -126 1119 -100
rect 1185 -122 1215 -100
rect 975 -172 991 -138
rect 1025 -172 1041 -138
rect 975 -188 1041 -172
rect 1167 -138 1233 -122
rect 1281 -126 1311 -100
rect 1377 -122 1407 -100
rect 1167 -172 1183 -138
rect 1217 -172 1233 -138
rect 1167 -188 1233 -172
rect 1359 -138 1425 -122
rect 1473 -126 1503 -100
rect 1569 -122 1599 -100
rect 1359 -172 1375 -138
rect 1409 -172 1425 -138
rect 1359 -188 1425 -172
rect 1551 -138 1617 -122
rect 1665 -126 1695 -100
rect 1761 -122 1791 -100
rect 1551 -172 1567 -138
rect 1601 -172 1617 -138
rect 1551 -188 1617 -172
rect 1743 -138 1809 -122
rect 1857 -126 1887 -100
rect 1953 -122 1983 -100
rect 1743 -172 1759 -138
rect 1793 -172 1809 -138
rect 1743 -188 1809 -172
rect 1935 -138 2001 -122
rect 2049 -126 2079 -100
rect 2145 -122 2175 -100
rect 1935 -172 1951 -138
rect 1985 -172 2001 -138
rect 1935 -188 2001 -172
rect 2127 -138 2193 -122
rect 2241 -126 2271 -100
rect 2337 -122 2367 -100
rect 2127 -172 2143 -138
rect 2177 -172 2193 -138
rect 2127 -188 2193 -172
rect 2319 -138 2385 -122
rect 2433 -126 2463 -100
rect 2529 -122 2559 -100
rect 2319 -172 2335 -138
rect 2369 -172 2385 -138
rect 2319 -188 2385 -172
rect 2511 -138 2577 -122
rect 2625 -126 2655 -100
rect 2721 -122 2751 -100
rect 2511 -172 2527 -138
rect 2561 -172 2577 -138
rect 2511 -188 2577 -172
rect 2703 -138 2769 -122
rect 2817 -126 2847 -100
rect 2703 -172 2719 -138
rect 2753 -172 2769 -138
rect 2703 -188 2769 -172
<< polycont >>
rect -2753 138 -2719 172
rect -2561 138 -2527 172
rect -2369 138 -2335 172
rect -2177 138 -2143 172
rect -1985 138 -1951 172
rect -1793 138 -1759 172
rect -1601 138 -1567 172
rect -1409 138 -1375 172
rect -1217 138 -1183 172
rect -1025 138 -991 172
rect -833 138 -799 172
rect -641 138 -607 172
rect -449 138 -415 172
rect -257 138 -223 172
rect -65 138 -31 172
rect 127 138 161 172
rect 319 138 353 172
rect 511 138 545 172
rect 703 138 737 172
rect 895 138 929 172
rect 1087 138 1121 172
rect 1279 138 1313 172
rect 1471 138 1505 172
rect 1663 138 1697 172
rect 1855 138 1889 172
rect 2047 138 2081 172
rect 2239 138 2273 172
rect 2431 138 2465 172
rect 2623 138 2657 172
rect 2815 138 2849 172
rect -2849 -172 -2815 -138
rect -2657 -172 -2623 -138
rect -2465 -172 -2431 -138
rect -2273 -172 -2239 -138
rect -2081 -172 -2047 -138
rect -1889 -172 -1855 -138
rect -1697 -172 -1663 -138
rect -1505 -172 -1471 -138
rect -1313 -172 -1279 -138
rect -1121 -172 -1087 -138
rect -929 -172 -895 -138
rect -737 -172 -703 -138
rect -545 -172 -511 -138
rect -353 -172 -319 -138
rect -161 -172 -127 -138
rect 31 -172 65 -138
rect 223 -172 257 -138
rect 415 -172 449 -138
rect 607 -172 641 -138
rect 799 -172 833 -138
rect 991 -172 1025 -138
rect 1183 -172 1217 -138
rect 1375 -172 1409 -138
rect 1567 -172 1601 -138
rect 1759 -172 1793 -138
rect 1951 -172 1985 -138
rect 2143 -172 2177 -138
rect 2335 -172 2369 -138
rect 2527 -172 2561 -138
rect 2719 -172 2753 -138
<< locali >>
rect -3011 240 -2915 274
rect 2915 240 3011 274
rect -3011 178 -2977 240
rect 2977 178 3011 240
rect -2769 138 -2753 172
rect -2719 138 -2703 172
rect -2577 138 -2561 172
rect -2527 138 -2511 172
rect -2385 138 -2369 172
rect -2335 138 -2319 172
rect -2193 138 -2177 172
rect -2143 138 -2127 172
rect -2001 138 -1985 172
rect -1951 138 -1935 172
rect -1809 138 -1793 172
rect -1759 138 -1743 172
rect -1617 138 -1601 172
rect -1567 138 -1551 172
rect -1425 138 -1409 172
rect -1375 138 -1359 172
rect -1233 138 -1217 172
rect -1183 138 -1167 172
rect -1041 138 -1025 172
rect -991 138 -975 172
rect -849 138 -833 172
rect -799 138 -783 172
rect -657 138 -641 172
rect -607 138 -591 172
rect -465 138 -449 172
rect -415 138 -399 172
rect -273 138 -257 172
rect -223 138 -207 172
rect -81 138 -65 172
rect -31 138 -15 172
rect 111 138 127 172
rect 161 138 177 172
rect 303 138 319 172
rect 353 138 369 172
rect 495 138 511 172
rect 545 138 561 172
rect 687 138 703 172
rect 737 138 753 172
rect 879 138 895 172
rect 929 138 945 172
rect 1071 138 1087 172
rect 1121 138 1137 172
rect 1263 138 1279 172
rect 1313 138 1329 172
rect 1455 138 1471 172
rect 1505 138 1521 172
rect 1647 138 1663 172
rect 1697 138 1713 172
rect 1839 138 1855 172
rect 1889 138 1905 172
rect 2031 138 2047 172
rect 2081 138 2097 172
rect 2223 138 2239 172
rect 2273 138 2289 172
rect 2415 138 2431 172
rect 2465 138 2481 172
rect 2607 138 2623 172
rect 2657 138 2673 172
rect 2799 138 2815 172
rect 2849 138 2865 172
rect -2897 88 -2863 104
rect -2897 -104 -2863 -88
rect -2801 88 -2767 104
rect -2801 -104 -2767 -88
rect -2705 88 -2671 104
rect -2705 -104 -2671 -88
rect -2609 88 -2575 104
rect -2609 -104 -2575 -88
rect -2513 88 -2479 104
rect -2513 -104 -2479 -88
rect -2417 88 -2383 104
rect -2417 -104 -2383 -88
rect -2321 88 -2287 104
rect -2321 -104 -2287 -88
rect -2225 88 -2191 104
rect -2225 -104 -2191 -88
rect -2129 88 -2095 104
rect -2129 -104 -2095 -88
rect -2033 88 -1999 104
rect -2033 -104 -1999 -88
rect -1937 88 -1903 104
rect -1937 -104 -1903 -88
rect -1841 88 -1807 104
rect -1841 -104 -1807 -88
rect -1745 88 -1711 104
rect -1745 -104 -1711 -88
rect -1649 88 -1615 104
rect -1649 -104 -1615 -88
rect -1553 88 -1519 104
rect -1553 -104 -1519 -88
rect -1457 88 -1423 104
rect -1457 -104 -1423 -88
rect -1361 88 -1327 104
rect -1361 -104 -1327 -88
rect -1265 88 -1231 104
rect -1265 -104 -1231 -88
rect -1169 88 -1135 104
rect -1169 -104 -1135 -88
rect -1073 88 -1039 104
rect -1073 -104 -1039 -88
rect -977 88 -943 104
rect -977 -104 -943 -88
rect -881 88 -847 104
rect -881 -104 -847 -88
rect -785 88 -751 104
rect -785 -104 -751 -88
rect -689 88 -655 104
rect -689 -104 -655 -88
rect -593 88 -559 104
rect -593 -104 -559 -88
rect -497 88 -463 104
rect -497 -104 -463 -88
rect -401 88 -367 104
rect -401 -104 -367 -88
rect -305 88 -271 104
rect -305 -104 -271 -88
rect -209 88 -175 104
rect -209 -104 -175 -88
rect -113 88 -79 104
rect -113 -104 -79 -88
rect -17 88 17 104
rect -17 -104 17 -88
rect 79 88 113 104
rect 79 -104 113 -88
rect 175 88 209 104
rect 175 -104 209 -88
rect 271 88 305 104
rect 271 -104 305 -88
rect 367 88 401 104
rect 367 -104 401 -88
rect 463 88 497 104
rect 463 -104 497 -88
rect 559 88 593 104
rect 559 -104 593 -88
rect 655 88 689 104
rect 655 -104 689 -88
rect 751 88 785 104
rect 751 -104 785 -88
rect 847 88 881 104
rect 847 -104 881 -88
rect 943 88 977 104
rect 943 -104 977 -88
rect 1039 88 1073 104
rect 1039 -104 1073 -88
rect 1135 88 1169 104
rect 1135 -104 1169 -88
rect 1231 88 1265 104
rect 1231 -104 1265 -88
rect 1327 88 1361 104
rect 1327 -104 1361 -88
rect 1423 88 1457 104
rect 1423 -104 1457 -88
rect 1519 88 1553 104
rect 1519 -104 1553 -88
rect 1615 88 1649 104
rect 1615 -104 1649 -88
rect 1711 88 1745 104
rect 1711 -104 1745 -88
rect 1807 88 1841 104
rect 1807 -104 1841 -88
rect 1903 88 1937 104
rect 1903 -104 1937 -88
rect 1999 88 2033 104
rect 1999 -104 2033 -88
rect 2095 88 2129 104
rect 2095 -104 2129 -88
rect 2191 88 2225 104
rect 2191 -104 2225 -88
rect 2287 88 2321 104
rect 2287 -104 2321 -88
rect 2383 88 2417 104
rect 2383 -104 2417 -88
rect 2479 88 2513 104
rect 2479 -104 2513 -88
rect 2575 88 2609 104
rect 2575 -104 2609 -88
rect 2671 88 2705 104
rect 2671 -104 2705 -88
rect 2767 88 2801 104
rect 2767 -104 2801 -88
rect 2863 88 2897 104
rect 2863 -104 2897 -88
rect -2865 -172 -2849 -138
rect -2815 -172 -2799 -138
rect -2673 -172 -2657 -138
rect -2623 -172 -2607 -138
rect -2481 -172 -2465 -138
rect -2431 -172 -2415 -138
rect -2289 -172 -2273 -138
rect -2239 -172 -2223 -138
rect -2097 -172 -2081 -138
rect -2047 -172 -2031 -138
rect -1905 -172 -1889 -138
rect -1855 -172 -1839 -138
rect -1713 -172 -1697 -138
rect -1663 -172 -1647 -138
rect -1521 -172 -1505 -138
rect -1471 -172 -1455 -138
rect -1329 -172 -1313 -138
rect -1279 -172 -1263 -138
rect -1137 -172 -1121 -138
rect -1087 -172 -1071 -138
rect -945 -172 -929 -138
rect -895 -172 -879 -138
rect -753 -172 -737 -138
rect -703 -172 -687 -138
rect -561 -172 -545 -138
rect -511 -172 -495 -138
rect -369 -172 -353 -138
rect -319 -172 -303 -138
rect -177 -172 -161 -138
rect -127 -172 -111 -138
rect 15 -172 31 -138
rect 65 -172 81 -138
rect 207 -172 223 -138
rect 257 -172 273 -138
rect 399 -172 415 -138
rect 449 -172 465 -138
rect 591 -172 607 -138
rect 641 -172 657 -138
rect 783 -172 799 -138
rect 833 -172 849 -138
rect 975 -172 991 -138
rect 1025 -172 1041 -138
rect 1167 -172 1183 -138
rect 1217 -172 1233 -138
rect 1359 -172 1375 -138
rect 1409 -172 1425 -138
rect 1551 -172 1567 -138
rect 1601 -172 1617 -138
rect 1743 -172 1759 -138
rect 1793 -172 1809 -138
rect 1935 -172 1951 -138
rect 1985 -172 2001 -138
rect 2127 -172 2143 -138
rect 2177 -172 2193 -138
rect 2319 -172 2335 -138
rect 2369 -172 2385 -138
rect 2511 -172 2527 -138
rect 2561 -172 2577 -138
rect 2703 -172 2719 -138
rect 2753 -172 2769 -138
rect -3011 -240 -2977 -178
rect 2977 -240 3011 -178
rect -3011 -274 -2915 -240
rect 2915 -274 3011 -240
<< viali >>
rect -2753 138 -2719 172
rect -2561 138 -2527 172
rect -2369 138 -2335 172
rect -2177 138 -2143 172
rect -1985 138 -1951 172
rect -1793 138 -1759 172
rect -1601 138 -1567 172
rect -1409 138 -1375 172
rect -1217 138 -1183 172
rect -1025 138 -991 172
rect -833 138 -799 172
rect -641 138 -607 172
rect -449 138 -415 172
rect -257 138 -223 172
rect -65 138 -31 172
rect 127 138 161 172
rect 319 138 353 172
rect 511 138 545 172
rect 703 138 737 172
rect 895 138 929 172
rect 1087 138 1121 172
rect 1279 138 1313 172
rect 1471 138 1505 172
rect 1663 138 1697 172
rect 1855 138 1889 172
rect 2047 138 2081 172
rect 2239 138 2273 172
rect 2431 138 2465 172
rect 2623 138 2657 172
rect 2815 138 2849 172
rect -2897 -88 -2863 88
rect -2801 -88 -2767 88
rect -2705 -88 -2671 88
rect -2609 -88 -2575 88
rect -2513 -88 -2479 88
rect -2417 -88 -2383 88
rect -2321 -88 -2287 88
rect -2225 -88 -2191 88
rect -2129 -88 -2095 88
rect -2033 -88 -1999 88
rect -1937 -88 -1903 88
rect -1841 -88 -1807 88
rect -1745 -88 -1711 88
rect -1649 -88 -1615 88
rect -1553 -88 -1519 88
rect -1457 -88 -1423 88
rect -1361 -88 -1327 88
rect -1265 -88 -1231 88
rect -1169 -88 -1135 88
rect -1073 -88 -1039 88
rect -977 -88 -943 88
rect -881 -88 -847 88
rect -785 -88 -751 88
rect -689 -88 -655 88
rect -593 -88 -559 88
rect -497 -88 -463 88
rect -401 -88 -367 88
rect -305 -88 -271 88
rect -209 -88 -175 88
rect -113 -88 -79 88
rect -17 -88 17 88
rect 79 -88 113 88
rect 175 -88 209 88
rect 271 -88 305 88
rect 367 -88 401 88
rect 463 -88 497 88
rect 559 -88 593 88
rect 655 -88 689 88
rect 751 -88 785 88
rect 847 -88 881 88
rect 943 -88 977 88
rect 1039 -88 1073 88
rect 1135 -88 1169 88
rect 1231 -88 1265 88
rect 1327 -88 1361 88
rect 1423 -88 1457 88
rect 1519 -88 1553 88
rect 1615 -88 1649 88
rect 1711 -88 1745 88
rect 1807 -88 1841 88
rect 1903 -88 1937 88
rect 1999 -88 2033 88
rect 2095 -88 2129 88
rect 2191 -88 2225 88
rect 2287 -88 2321 88
rect 2383 -88 2417 88
rect 2479 -88 2513 88
rect 2575 -88 2609 88
rect 2671 -88 2705 88
rect 2767 -88 2801 88
rect 2863 -88 2897 88
rect -2849 -172 -2815 -138
rect -2657 -172 -2623 -138
rect -2465 -172 -2431 -138
rect -2273 -172 -2239 -138
rect -2081 -172 -2047 -138
rect -1889 -172 -1855 -138
rect -1697 -172 -1663 -138
rect -1505 -172 -1471 -138
rect -1313 -172 -1279 -138
rect -1121 -172 -1087 -138
rect -929 -172 -895 -138
rect -737 -172 -703 -138
rect -545 -172 -511 -138
rect -353 -172 -319 -138
rect -161 -172 -127 -138
rect 31 -172 65 -138
rect 223 -172 257 -138
rect 415 -172 449 -138
rect 607 -172 641 -138
rect 799 -172 833 -138
rect 991 -172 1025 -138
rect 1183 -172 1217 -138
rect 1375 -172 1409 -138
rect 1567 -172 1601 -138
rect 1759 -172 1793 -138
rect 1951 -172 1985 -138
rect 2143 -172 2177 -138
rect 2335 -172 2369 -138
rect 2527 -172 2561 -138
rect 2719 -172 2753 -138
<< metal1 >>
rect -2765 172 -2707 178
rect -2765 138 -2753 172
rect -2719 138 -2707 172
rect -2765 132 -2707 138
rect -2573 172 -2515 178
rect -2573 138 -2561 172
rect -2527 138 -2515 172
rect -2573 132 -2515 138
rect -2381 172 -2323 178
rect -2381 138 -2369 172
rect -2335 138 -2323 172
rect -2381 132 -2323 138
rect -2189 172 -2131 178
rect -2189 138 -2177 172
rect -2143 138 -2131 172
rect -2189 132 -2131 138
rect -1997 172 -1939 178
rect -1997 138 -1985 172
rect -1951 138 -1939 172
rect -1997 132 -1939 138
rect -1805 172 -1747 178
rect -1805 138 -1793 172
rect -1759 138 -1747 172
rect -1805 132 -1747 138
rect -1613 172 -1555 178
rect -1613 138 -1601 172
rect -1567 138 -1555 172
rect -1613 132 -1555 138
rect -1421 172 -1363 178
rect -1421 138 -1409 172
rect -1375 138 -1363 172
rect -1421 132 -1363 138
rect -1229 172 -1171 178
rect -1229 138 -1217 172
rect -1183 138 -1171 172
rect -1229 132 -1171 138
rect -1037 172 -979 178
rect -1037 138 -1025 172
rect -991 138 -979 172
rect -1037 132 -979 138
rect -845 172 -787 178
rect -845 138 -833 172
rect -799 138 -787 172
rect -845 132 -787 138
rect -653 172 -595 178
rect -653 138 -641 172
rect -607 138 -595 172
rect -653 132 -595 138
rect -461 172 -403 178
rect -461 138 -449 172
rect -415 138 -403 172
rect -461 132 -403 138
rect -269 172 -211 178
rect -269 138 -257 172
rect -223 138 -211 172
rect -269 132 -211 138
rect -77 172 -19 178
rect -77 138 -65 172
rect -31 138 -19 172
rect -77 132 -19 138
rect 115 172 173 178
rect 115 138 127 172
rect 161 138 173 172
rect 115 132 173 138
rect 307 172 365 178
rect 307 138 319 172
rect 353 138 365 172
rect 307 132 365 138
rect 499 172 557 178
rect 499 138 511 172
rect 545 138 557 172
rect 499 132 557 138
rect 691 172 749 178
rect 691 138 703 172
rect 737 138 749 172
rect 691 132 749 138
rect 883 172 941 178
rect 883 138 895 172
rect 929 138 941 172
rect 883 132 941 138
rect 1075 172 1133 178
rect 1075 138 1087 172
rect 1121 138 1133 172
rect 1075 132 1133 138
rect 1267 172 1325 178
rect 1267 138 1279 172
rect 1313 138 1325 172
rect 1267 132 1325 138
rect 1459 172 1517 178
rect 1459 138 1471 172
rect 1505 138 1517 172
rect 1459 132 1517 138
rect 1651 172 1709 178
rect 1651 138 1663 172
rect 1697 138 1709 172
rect 1651 132 1709 138
rect 1843 172 1901 178
rect 1843 138 1855 172
rect 1889 138 1901 172
rect 1843 132 1901 138
rect 2035 172 2093 178
rect 2035 138 2047 172
rect 2081 138 2093 172
rect 2035 132 2093 138
rect 2227 172 2285 178
rect 2227 138 2239 172
rect 2273 138 2285 172
rect 2227 132 2285 138
rect 2419 172 2477 178
rect 2419 138 2431 172
rect 2465 138 2477 172
rect 2419 132 2477 138
rect 2611 172 2669 178
rect 2611 138 2623 172
rect 2657 138 2669 172
rect 2611 132 2669 138
rect 2803 172 2861 178
rect 2803 138 2815 172
rect 2849 138 2861 172
rect 2803 132 2861 138
rect -2903 88 -2857 100
rect -2903 -88 -2897 88
rect -2863 -88 -2857 88
rect -2903 -100 -2857 -88
rect -2807 88 -2761 100
rect -2807 -88 -2801 88
rect -2767 -88 -2761 88
rect -2807 -100 -2761 -88
rect -2711 88 -2665 100
rect -2711 -88 -2705 88
rect -2671 -88 -2665 88
rect -2711 -100 -2665 -88
rect -2615 88 -2569 100
rect -2615 -88 -2609 88
rect -2575 -88 -2569 88
rect -2615 -100 -2569 -88
rect -2519 88 -2473 100
rect -2519 -88 -2513 88
rect -2479 -88 -2473 88
rect -2519 -100 -2473 -88
rect -2423 88 -2377 100
rect -2423 -88 -2417 88
rect -2383 -88 -2377 88
rect -2423 -100 -2377 -88
rect -2327 88 -2281 100
rect -2327 -88 -2321 88
rect -2287 -88 -2281 88
rect -2327 -100 -2281 -88
rect -2231 88 -2185 100
rect -2231 -88 -2225 88
rect -2191 -88 -2185 88
rect -2231 -100 -2185 -88
rect -2135 88 -2089 100
rect -2135 -88 -2129 88
rect -2095 -88 -2089 88
rect -2135 -100 -2089 -88
rect -2039 88 -1993 100
rect -2039 -88 -2033 88
rect -1999 -88 -1993 88
rect -2039 -100 -1993 -88
rect -1943 88 -1897 100
rect -1943 -88 -1937 88
rect -1903 -88 -1897 88
rect -1943 -100 -1897 -88
rect -1847 88 -1801 100
rect -1847 -88 -1841 88
rect -1807 -88 -1801 88
rect -1847 -100 -1801 -88
rect -1751 88 -1705 100
rect -1751 -88 -1745 88
rect -1711 -88 -1705 88
rect -1751 -100 -1705 -88
rect -1655 88 -1609 100
rect -1655 -88 -1649 88
rect -1615 -88 -1609 88
rect -1655 -100 -1609 -88
rect -1559 88 -1513 100
rect -1559 -88 -1553 88
rect -1519 -88 -1513 88
rect -1559 -100 -1513 -88
rect -1463 88 -1417 100
rect -1463 -88 -1457 88
rect -1423 -88 -1417 88
rect -1463 -100 -1417 -88
rect -1367 88 -1321 100
rect -1367 -88 -1361 88
rect -1327 -88 -1321 88
rect -1367 -100 -1321 -88
rect -1271 88 -1225 100
rect -1271 -88 -1265 88
rect -1231 -88 -1225 88
rect -1271 -100 -1225 -88
rect -1175 88 -1129 100
rect -1175 -88 -1169 88
rect -1135 -88 -1129 88
rect -1175 -100 -1129 -88
rect -1079 88 -1033 100
rect -1079 -88 -1073 88
rect -1039 -88 -1033 88
rect -1079 -100 -1033 -88
rect -983 88 -937 100
rect -983 -88 -977 88
rect -943 -88 -937 88
rect -983 -100 -937 -88
rect -887 88 -841 100
rect -887 -88 -881 88
rect -847 -88 -841 88
rect -887 -100 -841 -88
rect -791 88 -745 100
rect -791 -88 -785 88
rect -751 -88 -745 88
rect -791 -100 -745 -88
rect -695 88 -649 100
rect -695 -88 -689 88
rect -655 -88 -649 88
rect -695 -100 -649 -88
rect -599 88 -553 100
rect -599 -88 -593 88
rect -559 -88 -553 88
rect -599 -100 -553 -88
rect -503 88 -457 100
rect -503 -88 -497 88
rect -463 -88 -457 88
rect -503 -100 -457 -88
rect -407 88 -361 100
rect -407 -88 -401 88
rect -367 -88 -361 88
rect -407 -100 -361 -88
rect -311 88 -265 100
rect -311 -88 -305 88
rect -271 -88 -265 88
rect -311 -100 -265 -88
rect -215 88 -169 100
rect -215 -88 -209 88
rect -175 -88 -169 88
rect -215 -100 -169 -88
rect -119 88 -73 100
rect -119 -88 -113 88
rect -79 -88 -73 88
rect -119 -100 -73 -88
rect -23 88 23 100
rect -23 -88 -17 88
rect 17 -88 23 88
rect -23 -100 23 -88
rect 73 88 119 100
rect 73 -88 79 88
rect 113 -88 119 88
rect 73 -100 119 -88
rect 169 88 215 100
rect 169 -88 175 88
rect 209 -88 215 88
rect 169 -100 215 -88
rect 265 88 311 100
rect 265 -88 271 88
rect 305 -88 311 88
rect 265 -100 311 -88
rect 361 88 407 100
rect 361 -88 367 88
rect 401 -88 407 88
rect 361 -100 407 -88
rect 457 88 503 100
rect 457 -88 463 88
rect 497 -88 503 88
rect 457 -100 503 -88
rect 553 88 599 100
rect 553 -88 559 88
rect 593 -88 599 88
rect 553 -100 599 -88
rect 649 88 695 100
rect 649 -88 655 88
rect 689 -88 695 88
rect 649 -100 695 -88
rect 745 88 791 100
rect 745 -88 751 88
rect 785 -88 791 88
rect 745 -100 791 -88
rect 841 88 887 100
rect 841 -88 847 88
rect 881 -88 887 88
rect 841 -100 887 -88
rect 937 88 983 100
rect 937 -88 943 88
rect 977 -88 983 88
rect 937 -100 983 -88
rect 1033 88 1079 100
rect 1033 -88 1039 88
rect 1073 -88 1079 88
rect 1033 -100 1079 -88
rect 1129 88 1175 100
rect 1129 -88 1135 88
rect 1169 -88 1175 88
rect 1129 -100 1175 -88
rect 1225 88 1271 100
rect 1225 -88 1231 88
rect 1265 -88 1271 88
rect 1225 -100 1271 -88
rect 1321 88 1367 100
rect 1321 -88 1327 88
rect 1361 -88 1367 88
rect 1321 -100 1367 -88
rect 1417 88 1463 100
rect 1417 -88 1423 88
rect 1457 -88 1463 88
rect 1417 -100 1463 -88
rect 1513 88 1559 100
rect 1513 -88 1519 88
rect 1553 -88 1559 88
rect 1513 -100 1559 -88
rect 1609 88 1655 100
rect 1609 -88 1615 88
rect 1649 -88 1655 88
rect 1609 -100 1655 -88
rect 1705 88 1751 100
rect 1705 -88 1711 88
rect 1745 -88 1751 88
rect 1705 -100 1751 -88
rect 1801 88 1847 100
rect 1801 -88 1807 88
rect 1841 -88 1847 88
rect 1801 -100 1847 -88
rect 1897 88 1943 100
rect 1897 -88 1903 88
rect 1937 -88 1943 88
rect 1897 -100 1943 -88
rect 1993 88 2039 100
rect 1993 -88 1999 88
rect 2033 -88 2039 88
rect 1993 -100 2039 -88
rect 2089 88 2135 100
rect 2089 -88 2095 88
rect 2129 -88 2135 88
rect 2089 -100 2135 -88
rect 2185 88 2231 100
rect 2185 -88 2191 88
rect 2225 -88 2231 88
rect 2185 -100 2231 -88
rect 2281 88 2327 100
rect 2281 -88 2287 88
rect 2321 -88 2327 88
rect 2281 -100 2327 -88
rect 2377 88 2423 100
rect 2377 -88 2383 88
rect 2417 -88 2423 88
rect 2377 -100 2423 -88
rect 2473 88 2519 100
rect 2473 -88 2479 88
rect 2513 -88 2519 88
rect 2473 -100 2519 -88
rect 2569 88 2615 100
rect 2569 -88 2575 88
rect 2609 -88 2615 88
rect 2569 -100 2615 -88
rect 2665 88 2711 100
rect 2665 -88 2671 88
rect 2705 -88 2711 88
rect 2665 -100 2711 -88
rect 2761 88 2807 100
rect 2761 -88 2767 88
rect 2801 -88 2807 88
rect 2761 -100 2807 -88
rect 2857 88 2903 100
rect 2857 -88 2863 88
rect 2897 -88 2903 88
rect 2857 -100 2903 -88
rect -2861 -138 -2803 -132
rect -2861 -172 -2849 -138
rect -2815 -172 -2803 -138
rect -2861 -178 -2803 -172
rect -2669 -138 -2611 -132
rect -2669 -172 -2657 -138
rect -2623 -172 -2611 -138
rect -2669 -178 -2611 -172
rect -2477 -138 -2419 -132
rect -2477 -172 -2465 -138
rect -2431 -172 -2419 -138
rect -2477 -178 -2419 -172
rect -2285 -138 -2227 -132
rect -2285 -172 -2273 -138
rect -2239 -172 -2227 -138
rect -2285 -178 -2227 -172
rect -2093 -138 -2035 -132
rect -2093 -172 -2081 -138
rect -2047 -172 -2035 -138
rect -2093 -178 -2035 -172
rect -1901 -138 -1843 -132
rect -1901 -172 -1889 -138
rect -1855 -172 -1843 -138
rect -1901 -178 -1843 -172
rect -1709 -138 -1651 -132
rect -1709 -172 -1697 -138
rect -1663 -172 -1651 -138
rect -1709 -178 -1651 -172
rect -1517 -138 -1459 -132
rect -1517 -172 -1505 -138
rect -1471 -172 -1459 -138
rect -1517 -178 -1459 -172
rect -1325 -138 -1267 -132
rect -1325 -172 -1313 -138
rect -1279 -172 -1267 -138
rect -1325 -178 -1267 -172
rect -1133 -138 -1075 -132
rect -1133 -172 -1121 -138
rect -1087 -172 -1075 -138
rect -1133 -178 -1075 -172
rect -941 -138 -883 -132
rect -941 -172 -929 -138
rect -895 -172 -883 -138
rect -941 -178 -883 -172
rect -749 -138 -691 -132
rect -749 -172 -737 -138
rect -703 -172 -691 -138
rect -749 -178 -691 -172
rect -557 -138 -499 -132
rect -557 -172 -545 -138
rect -511 -172 -499 -138
rect -557 -178 -499 -172
rect -365 -138 -307 -132
rect -365 -172 -353 -138
rect -319 -172 -307 -138
rect -365 -178 -307 -172
rect -173 -138 -115 -132
rect -173 -172 -161 -138
rect -127 -172 -115 -138
rect -173 -178 -115 -172
rect 19 -138 77 -132
rect 19 -172 31 -138
rect 65 -172 77 -138
rect 19 -178 77 -172
rect 211 -138 269 -132
rect 211 -172 223 -138
rect 257 -172 269 -138
rect 211 -178 269 -172
rect 403 -138 461 -132
rect 403 -172 415 -138
rect 449 -172 461 -138
rect 403 -178 461 -172
rect 595 -138 653 -132
rect 595 -172 607 -138
rect 641 -172 653 -138
rect 595 -178 653 -172
rect 787 -138 845 -132
rect 787 -172 799 -138
rect 833 -172 845 -138
rect 787 -178 845 -172
rect 979 -138 1037 -132
rect 979 -172 991 -138
rect 1025 -172 1037 -138
rect 979 -178 1037 -172
rect 1171 -138 1229 -132
rect 1171 -172 1183 -138
rect 1217 -172 1229 -138
rect 1171 -178 1229 -172
rect 1363 -138 1421 -132
rect 1363 -172 1375 -138
rect 1409 -172 1421 -138
rect 1363 -178 1421 -172
rect 1555 -138 1613 -132
rect 1555 -172 1567 -138
rect 1601 -172 1613 -138
rect 1555 -178 1613 -172
rect 1747 -138 1805 -132
rect 1747 -172 1759 -138
rect 1793 -172 1805 -138
rect 1747 -178 1805 -172
rect 1939 -138 1997 -132
rect 1939 -172 1951 -138
rect 1985 -172 1997 -138
rect 1939 -178 1997 -172
rect 2131 -138 2189 -132
rect 2131 -172 2143 -138
rect 2177 -172 2189 -138
rect 2131 -178 2189 -172
rect 2323 -138 2381 -132
rect 2323 -172 2335 -138
rect 2369 -172 2381 -138
rect 2323 -178 2381 -172
rect 2515 -138 2573 -132
rect 2515 -172 2527 -138
rect 2561 -172 2573 -138
rect 2515 -178 2573 -172
rect 2707 -138 2765 -132
rect 2707 -172 2719 -138
rect 2753 -172 2765 -138
rect 2707 -178 2765 -172
<< properties >>
string FIXED_BBOX -2994 -257 2994 257
string gencell sky130_fd_pr__nfet_01v8_lvt
string library sky130
string parameters w 1.0 l 0.15 m 1 nf 60 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
