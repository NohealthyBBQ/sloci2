magic
tech sky130A
timestamp 1672463399
<< pwell >>
rect -325 -325 325 325
<< psubdiff >>
rect -307 301 307 307
rect -307 284 -253 301
rect 253 284 307 301
rect -307 278 307 284
rect -307 253 -278 278
rect -307 -253 -301 253
rect -284 -253 -278 253
rect 278 253 307 278
rect -307 -278 -278 -253
rect 278 -253 284 253
rect 301 -253 307 253
rect 278 -278 307 -253
rect -307 -284 307 -278
rect -307 -301 -253 -284
rect 253 -301 307 -284
rect -307 -307 307 -301
<< psubdiffcont >>
rect -253 284 253 301
rect -301 -253 -284 253
rect 284 -253 301 253
rect -253 -301 253 -284
<< ndiodelvt >>
rect -250 244 250 250
rect -250 -244 -244 244
rect 244 -244 250 244
rect -250 -250 250 -244
<< ndiodelvtc >>
rect -244 -244 244 244
<< locali >>
rect -301 284 -253 301
rect 253 284 301 301
rect -301 253 -284 284
rect 284 253 301 284
rect -252 -244 -244 244
rect 244 -244 252 244
rect -301 -284 -284 -253
rect 284 -284 301 -253
rect -301 -301 -253 -284
rect 253 -301 301 -284
<< viali >>
rect -244 -244 244 244
<< metal1 >>
rect -250 244 250 247
rect -250 -244 -244 244
rect 244 -244 250 244
rect -250 -247 250 -244
<< properties >>
string FIXED_BBOX -292 -292 292 292
string gencell sky130_fd_pr__diode_pw2nd_05v5_lvt
string library sky130
string parameters w 5 l 5 area 25.0 peri 20.0 nx 1 ny 1 dummy 0 lmin 0.45 wmin 0.45 elc 1 erc 1 etc 1 ebc 1 doverlap 0 compatible {sky130_fd_pr__diode_pw2nd_05v5 sky130_fd_pr__diode_pw2nd_05v5_lvt  sky130_fd_pr__diode_pw2nd_05v5_nvt sky130_fd_pr__diode_pw2nd_11v0} full_metal 1 vias 1 viagb 0 viagt 0 viagl 0 viagr 0
<< end >>
