magic
tech sky130A
magscale 1 2
timestamp 1662404926
<< error_p >>
rect -927 181 -865 187
rect -799 181 -737 187
rect -671 181 -609 187
rect -543 181 -481 187
rect -415 181 -353 187
rect -287 181 -225 187
rect -159 181 -97 187
rect -31 181 31 187
rect 97 181 159 187
rect 225 181 287 187
rect 353 181 415 187
rect 481 181 543 187
rect 609 181 671 187
rect 737 181 799 187
rect 865 181 927 187
rect -927 147 -915 181
rect -799 147 -787 181
rect -671 147 -659 181
rect -543 147 -531 181
rect -415 147 -403 181
rect -287 147 -275 181
rect -159 147 -147 181
rect -31 147 -19 181
rect 97 147 109 181
rect 225 147 237 181
rect 353 147 365 181
rect 481 147 493 181
rect 609 147 621 181
rect 737 147 749 181
rect 865 147 877 181
rect -927 141 -865 147
rect -799 141 -737 147
rect -671 141 -609 147
rect -543 141 -481 147
rect -415 141 -353 147
rect -287 141 -225 147
rect -159 141 -97 147
rect -31 141 31 147
rect 97 141 159 147
rect 225 141 287 147
rect 353 141 415 147
rect 481 141 543 147
rect 609 141 671 147
rect 737 141 799 147
rect 865 141 927 147
rect -927 -147 -865 -141
rect -799 -147 -737 -141
rect -671 -147 -609 -141
rect -543 -147 -481 -141
rect -415 -147 -353 -141
rect -287 -147 -225 -141
rect -159 -147 -97 -141
rect -31 -147 31 -141
rect 97 -147 159 -141
rect 225 -147 287 -141
rect 353 -147 415 -141
rect 481 -147 543 -141
rect 609 -147 671 -141
rect 737 -147 799 -141
rect 865 -147 927 -141
rect -927 -181 -915 -147
rect -799 -181 -787 -147
rect -671 -181 -659 -147
rect -543 -181 -531 -147
rect -415 -181 -403 -147
rect -287 -181 -275 -147
rect -159 -181 -147 -147
rect -31 -181 -19 -147
rect 97 -181 109 -147
rect 225 -181 237 -147
rect 353 -181 365 -147
rect 481 -181 493 -147
rect 609 -181 621 -147
rect 737 -181 749 -147
rect 865 -181 877 -147
rect -927 -187 -865 -181
rect -799 -187 -737 -181
rect -671 -187 -609 -181
rect -543 -187 -481 -181
rect -415 -187 -353 -181
rect -287 -187 -225 -181
rect -159 -187 -97 -181
rect -31 -187 31 -181
rect 97 -187 159 -181
rect 225 -187 287 -181
rect 353 -187 415 -181
rect 481 -187 543 -181
rect 609 -187 671 -181
rect 737 -187 799 -181
rect 865 -187 927 -181
<< nwell >>
rect -1127 -319 1127 319
<< pmoslvt >>
rect -931 -100 -861 100
rect -803 -100 -733 100
rect -675 -100 -605 100
rect -547 -100 -477 100
rect -419 -100 -349 100
rect -291 -100 -221 100
rect -163 -100 -93 100
rect -35 -100 35 100
rect 93 -100 163 100
rect 221 -100 291 100
rect 349 -100 419 100
rect 477 -100 547 100
rect 605 -100 675 100
rect 733 -100 803 100
rect 861 -100 931 100
<< pdiff >>
rect -989 88 -931 100
rect -989 -88 -977 88
rect -943 -88 -931 88
rect -989 -100 -931 -88
rect -861 88 -803 100
rect -861 -88 -849 88
rect -815 -88 -803 88
rect -861 -100 -803 -88
rect -733 88 -675 100
rect -733 -88 -721 88
rect -687 -88 -675 88
rect -733 -100 -675 -88
rect -605 88 -547 100
rect -605 -88 -593 88
rect -559 -88 -547 88
rect -605 -100 -547 -88
rect -477 88 -419 100
rect -477 -88 -465 88
rect -431 -88 -419 88
rect -477 -100 -419 -88
rect -349 88 -291 100
rect -349 -88 -337 88
rect -303 -88 -291 88
rect -349 -100 -291 -88
rect -221 88 -163 100
rect -221 -88 -209 88
rect -175 -88 -163 88
rect -221 -100 -163 -88
rect -93 88 -35 100
rect -93 -88 -81 88
rect -47 -88 -35 88
rect -93 -100 -35 -88
rect 35 88 93 100
rect 35 -88 47 88
rect 81 -88 93 88
rect 35 -100 93 -88
rect 163 88 221 100
rect 163 -88 175 88
rect 209 -88 221 88
rect 163 -100 221 -88
rect 291 88 349 100
rect 291 -88 303 88
rect 337 -88 349 88
rect 291 -100 349 -88
rect 419 88 477 100
rect 419 -88 431 88
rect 465 -88 477 88
rect 419 -100 477 -88
rect 547 88 605 100
rect 547 -88 559 88
rect 593 -88 605 88
rect 547 -100 605 -88
rect 675 88 733 100
rect 675 -88 687 88
rect 721 -88 733 88
rect 675 -100 733 -88
rect 803 88 861 100
rect 803 -88 815 88
rect 849 -88 861 88
rect 803 -100 861 -88
rect 931 88 989 100
rect 931 -88 943 88
rect 977 -88 989 88
rect 931 -100 989 -88
<< pdiffc >>
rect -977 -88 -943 88
rect -849 -88 -815 88
rect -721 -88 -687 88
rect -593 -88 -559 88
rect -465 -88 -431 88
rect -337 -88 -303 88
rect -209 -88 -175 88
rect -81 -88 -47 88
rect 47 -88 81 88
rect 175 -88 209 88
rect 303 -88 337 88
rect 431 -88 465 88
rect 559 -88 593 88
rect 687 -88 721 88
rect 815 -88 849 88
rect 943 -88 977 88
<< nsubdiff >>
rect -1091 249 -995 283
rect 995 249 1091 283
rect -1091 187 -1057 249
rect 1057 187 1091 249
rect -1091 -249 -1057 -187
rect 1057 -249 1091 -187
rect -1091 -283 -995 -249
rect 995 -283 1091 -249
<< nsubdiffcont >>
rect -995 249 995 283
rect -1091 -187 -1057 187
rect 1057 -187 1091 187
rect -995 -283 995 -249
<< poly >>
rect -931 181 -861 197
rect -931 147 -915 181
rect -877 147 -861 181
rect -931 100 -861 147
rect -803 181 -733 197
rect -803 147 -787 181
rect -749 147 -733 181
rect -803 100 -733 147
rect -675 181 -605 197
rect -675 147 -659 181
rect -621 147 -605 181
rect -675 100 -605 147
rect -547 181 -477 197
rect -547 147 -531 181
rect -493 147 -477 181
rect -547 100 -477 147
rect -419 181 -349 197
rect -419 147 -403 181
rect -365 147 -349 181
rect -419 100 -349 147
rect -291 181 -221 197
rect -291 147 -275 181
rect -237 147 -221 181
rect -291 100 -221 147
rect -163 181 -93 197
rect -163 147 -147 181
rect -109 147 -93 181
rect -163 100 -93 147
rect -35 181 35 197
rect -35 147 -19 181
rect 19 147 35 181
rect -35 100 35 147
rect 93 181 163 197
rect 93 147 109 181
rect 147 147 163 181
rect 93 100 163 147
rect 221 181 291 197
rect 221 147 237 181
rect 275 147 291 181
rect 221 100 291 147
rect 349 181 419 197
rect 349 147 365 181
rect 403 147 419 181
rect 349 100 419 147
rect 477 181 547 197
rect 477 147 493 181
rect 531 147 547 181
rect 477 100 547 147
rect 605 181 675 197
rect 605 147 621 181
rect 659 147 675 181
rect 605 100 675 147
rect 733 181 803 197
rect 733 147 749 181
rect 787 147 803 181
rect 733 100 803 147
rect 861 181 931 197
rect 861 147 877 181
rect 915 147 931 181
rect 861 100 931 147
rect -931 -147 -861 -100
rect -931 -181 -915 -147
rect -877 -181 -861 -147
rect -931 -197 -861 -181
rect -803 -147 -733 -100
rect -803 -181 -787 -147
rect -749 -181 -733 -147
rect -803 -197 -733 -181
rect -675 -147 -605 -100
rect -675 -181 -659 -147
rect -621 -181 -605 -147
rect -675 -197 -605 -181
rect -547 -147 -477 -100
rect -547 -181 -531 -147
rect -493 -181 -477 -147
rect -547 -197 -477 -181
rect -419 -147 -349 -100
rect -419 -181 -403 -147
rect -365 -181 -349 -147
rect -419 -197 -349 -181
rect -291 -147 -221 -100
rect -291 -181 -275 -147
rect -237 -181 -221 -147
rect -291 -197 -221 -181
rect -163 -147 -93 -100
rect -163 -181 -147 -147
rect -109 -181 -93 -147
rect -163 -197 -93 -181
rect -35 -147 35 -100
rect -35 -181 -19 -147
rect 19 -181 35 -147
rect -35 -197 35 -181
rect 93 -147 163 -100
rect 93 -181 109 -147
rect 147 -181 163 -147
rect 93 -197 163 -181
rect 221 -147 291 -100
rect 221 -181 237 -147
rect 275 -181 291 -147
rect 221 -197 291 -181
rect 349 -147 419 -100
rect 349 -181 365 -147
rect 403 -181 419 -147
rect 349 -197 419 -181
rect 477 -147 547 -100
rect 477 -181 493 -147
rect 531 -181 547 -147
rect 477 -197 547 -181
rect 605 -147 675 -100
rect 605 -181 621 -147
rect 659 -181 675 -147
rect 605 -197 675 -181
rect 733 -147 803 -100
rect 733 -181 749 -147
rect 787 -181 803 -147
rect 733 -197 803 -181
rect 861 -147 931 -100
rect 861 -181 877 -147
rect 915 -181 931 -147
rect 861 -197 931 -181
<< polycont >>
rect -915 147 -877 181
rect -787 147 -749 181
rect -659 147 -621 181
rect -531 147 -493 181
rect -403 147 -365 181
rect -275 147 -237 181
rect -147 147 -109 181
rect -19 147 19 181
rect 109 147 147 181
rect 237 147 275 181
rect 365 147 403 181
rect 493 147 531 181
rect 621 147 659 181
rect 749 147 787 181
rect 877 147 915 181
rect -915 -181 -877 -147
rect -787 -181 -749 -147
rect -659 -181 -621 -147
rect -531 -181 -493 -147
rect -403 -181 -365 -147
rect -275 -181 -237 -147
rect -147 -181 -109 -147
rect -19 -181 19 -147
rect 109 -181 147 -147
rect 237 -181 275 -147
rect 365 -181 403 -147
rect 493 -181 531 -147
rect 621 -181 659 -147
rect 749 -181 787 -147
rect 877 -181 915 -147
<< locali >>
rect -1091 249 -995 283
rect 995 249 1091 283
rect -1091 187 -1057 249
rect 1057 187 1091 249
rect -931 147 -915 181
rect -877 147 -861 181
rect -803 147 -787 181
rect -749 147 -733 181
rect -675 147 -659 181
rect -621 147 -605 181
rect -547 147 -531 181
rect -493 147 -477 181
rect -419 147 -403 181
rect -365 147 -349 181
rect -291 147 -275 181
rect -237 147 -221 181
rect -163 147 -147 181
rect -109 147 -93 181
rect -35 147 -19 181
rect 19 147 35 181
rect 93 147 109 181
rect 147 147 163 181
rect 221 147 237 181
rect 275 147 291 181
rect 349 147 365 181
rect 403 147 419 181
rect 477 147 493 181
rect 531 147 547 181
rect 605 147 621 181
rect 659 147 675 181
rect 733 147 749 181
rect 787 147 803 181
rect 861 147 877 181
rect 915 147 931 181
rect -977 88 -943 104
rect -977 -104 -943 -88
rect -849 88 -815 104
rect -849 -104 -815 -88
rect -721 88 -687 104
rect -721 -104 -687 -88
rect -593 88 -559 104
rect -593 -104 -559 -88
rect -465 88 -431 104
rect -465 -104 -431 -88
rect -337 88 -303 104
rect -337 -104 -303 -88
rect -209 88 -175 104
rect -209 -104 -175 -88
rect -81 88 -47 104
rect -81 -104 -47 -88
rect 47 88 81 104
rect 47 -104 81 -88
rect 175 88 209 104
rect 175 -104 209 -88
rect 303 88 337 104
rect 303 -104 337 -88
rect 431 88 465 104
rect 431 -104 465 -88
rect 559 88 593 104
rect 559 -104 593 -88
rect 687 88 721 104
rect 687 -104 721 -88
rect 815 88 849 104
rect 815 -104 849 -88
rect 943 88 977 104
rect 943 -104 977 -88
rect -931 -181 -915 -147
rect -877 -181 -861 -147
rect -803 -181 -787 -147
rect -749 -181 -733 -147
rect -675 -181 -659 -147
rect -621 -181 -605 -147
rect -547 -181 -531 -147
rect -493 -181 -477 -147
rect -419 -181 -403 -147
rect -365 -181 -349 -147
rect -291 -181 -275 -147
rect -237 -181 -221 -147
rect -163 -181 -147 -147
rect -109 -181 -93 -147
rect -35 -181 -19 -147
rect 19 -181 35 -147
rect 93 -181 109 -147
rect 147 -181 163 -147
rect 221 -181 237 -147
rect 275 -181 291 -147
rect 349 -181 365 -147
rect 403 -181 419 -147
rect 477 -181 493 -147
rect 531 -181 547 -147
rect 605 -181 621 -147
rect 659 -181 675 -147
rect 733 -181 749 -147
rect 787 -181 803 -147
rect 861 -181 877 -147
rect 915 -181 931 -147
rect -1091 -249 -1057 -187
rect 1057 -249 1091 -187
rect -1091 -283 -995 -249
rect 995 -283 1091 -249
<< viali >>
rect -915 147 -877 181
rect -787 147 -749 181
rect -659 147 -621 181
rect -531 147 -493 181
rect -403 147 -365 181
rect -275 147 -237 181
rect -147 147 -109 181
rect -19 147 19 181
rect 109 147 147 181
rect 237 147 275 181
rect 365 147 403 181
rect 493 147 531 181
rect 621 147 659 181
rect 749 147 787 181
rect 877 147 915 181
rect -977 -88 -943 88
rect -849 -88 -815 88
rect -721 -88 -687 88
rect -593 -88 -559 88
rect -465 -88 -431 88
rect -337 -88 -303 88
rect -209 -88 -175 88
rect -81 -88 -47 88
rect 47 -88 81 88
rect 175 -88 209 88
rect 303 -88 337 88
rect 431 -88 465 88
rect 559 -88 593 88
rect 687 -88 721 88
rect 815 -88 849 88
rect 943 -88 977 88
rect -915 -181 -877 -147
rect -787 -181 -749 -147
rect -659 -181 -621 -147
rect -531 -181 -493 -147
rect -403 -181 -365 -147
rect -275 -181 -237 -147
rect -147 -181 -109 -147
rect -19 -181 19 -147
rect 109 -181 147 -147
rect 237 -181 275 -147
rect 365 -181 403 -147
rect 493 -181 531 -147
rect 621 -181 659 -147
rect 749 -181 787 -147
rect 877 -181 915 -147
<< metal1 >>
rect -927 181 -865 187
rect -927 147 -915 181
rect -877 147 -865 181
rect -927 141 -865 147
rect -799 181 -737 187
rect -799 147 -787 181
rect -749 147 -737 181
rect -799 141 -737 147
rect -671 181 -609 187
rect -671 147 -659 181
rect -621 147 -609 181
rect -671 141 -609 147
rect -543 181 -481 187
rect -543 147 -531 181
rect -493 147 -481 181
rect -543 141 -481 147
rect -415 181 -353 187
rect -415 147 -403 181
rect -365 147 -353 181
rect -415 141 -353 147
rect -287 181 -225 187
rect -287 147 -275 181
rect -237 147 -225 181
rect -287 141 -225 147
rect -159 181 -97 187
rect -159 147 -147 181
rect -109 147 -97 181
rect -159 141 -97 147
rect -31 181 31 187
rect -31 147 -19 181
rect 19 147 31 181
rect -31 141 31 147
rect 97 181 159 187
rect 97 147 109 181
rect 147 147 159 181
rect 97 141 159 147
rect 225 181 287 187
rect 225 147 237 181
rect 275 147 287 181
rect 225 141 287 147
rect 353 181 415 187
rect 353 147 365 181
rect 403 147 415 181
rect 353 141 415 147
rect 481 181 543 187
rect 481 147 493 181
rect 531 147 543 181
rect 481 141 543 147
rect 609 181 671 187
rect 609 147 621 181
rect 659 147 671 181
rect 609 141 671 147
rect 737 181 799 187
rect 737 147 749 181
rect 787 147 799 181
rect 737 141 799 147
rect 865 181 927 187
rect 865 147 877 181
rect 915 147 927 181
rect 865 141 927 147
rect -983 88 -937 100
rect -983 -88 -977 88
rect -943 -88 -937 88
rect -983 -100 -937 -88
rect -855 88 -809 100
rect -855 -88 -849 88
rect -815 -88 -809 88
rect -855 -100 -809 -88
rect -727 88 -681 100
rect -727 -88 -721 88
rect -687 -88 -681 88
rect -727 -100 -681 -88
rect -599 88 -553 100
rect -599 -88 -593 88
rect -559 -88 -553 88
rect -599 -100 -553 -88
rect -471 88 -425 100
rect -471 -88 -465 88
rect -431 -88 -425 88
rect -471 -100 -425 -88
rect -343 88 -297 100
rect -343 -88 -337 88
rect -303 -88 -297 88
rect -343 -100 -297 -88
rect -215 88 -169 100
rect -215 -88 -209 88
rect -175 -88 -169 88
rect -215 -100 -169 -88
rect -87 88 -41 100
rect -87 -88 -81 88
rect -47 -88 -41 88
rect -87 -100 -41 -88
rect 41 88 87 100
rect 41 -88 47 88
rect 81 -88 87 88
rect 41 -100 87 -88
rect 169 88 215 100
rect 169 -88 175 88
rect 209 -88 215 88
rect 169 -100 215 -88
rect 297 88 343 100
rect 297 -88 303 88
rect 337 -88 343 88
rect 297 -100 343 -88
rect 425 88 471 100
rect 425 -88 431 88
rect 465 -88 471 88
rect 425 -100 471 -88
rect 553 88 599 100
rect 553 -88 559 88
rect 593 -88 599 88
rect 553 -100 599 -88
rect 681 88 727 100
rect 681 -88 687 88
rect 721 -88 727 88
rect 681 -100 727 -88
rect 809 88 855 100
rect 809 -88 815 88
rect 849 -88 855 88
rect 809 -100 855 -88
rect 937 88 983 100
rect 937 -88 943 88
rect 977 -88 983 88
rect 937 -100 983 -88
rect -927 -147 -865 -141
rect -927 -181 -915 -147
rect -877 -181 -865 -147
rect -927 -187 -865 -181
rect -799 -147 -737 -141
rect -799 -181 -787 -147
rect -749 -181 -737 -147
rect -799 -187 -737 -181
rect -671 -147 -609 -141
rect -671 -181 -659 -147
rect -621 -181 -609 -147
rect -671 -187 -609 -181
rect -543 -147 -481 -141
rect -543 -181 -531 -147
rect -493 -181 -481 -147
rect -543 -187 -481 -181
rect -415 -147 -353 -141
rect -415 -181 -403 -147
rect -365 -181 -353 -147
rect -415 -187 -353 -181
rect -287 -147 -225 -141
rect -287 -181 -275 -147
rect -237 -181 -225 -147
rect -287 -187 -225 -181
rect -159 -147 -97 -141
rect -159 -181 -147 -147
rect -109 -181 -97 -147
rect -159 -187 -97 -181
rect -31 -147 31 -141
rect -31 -181 -19 -147
rect 19 -181 31 -147
rect -31 -187 31 -181
rect 97 -147 159 -141
rect 97 -181 109 -147
rect 147 -181 159 -147
rect 97 -187 159 -181
rect 225 -147 287 -141
rect 225 -181 237 -147
rect 275 -181 287 -147
rect 225 -187 287 -181
rect 353 -147 415 -141
rect 353 -181 365 -147
rect 403 -181 415 -147
rect 353 -187 415 -181
rect 481 -147 543 -141
rect 481 -181 493 -147
rect 531 -181 543 -147
rect 481 -187 543 -181
rect 609 -147 671 -141
rect 609 -181 621 -147
rect 659 -181 671 -147
rect 609 -187 671 -181
rect 737 -147 799 -141
rect 737 -181 749 -147
rect 787 -181 799 -147
rect 737 -187 799 -181
rect 865 -147 927 -141
rect 865 -181 877 -147
rect 915 -181 927 -147
rect 865 -187 927 -181
<< properties >>
string FIXED_BBOX -1074 -266 1074 266
string gencell sky130_fd_pr__pfet_01v8_lvt
string library sky130
string parameters w 1.0 l 0.35 m 1 nf 15 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.35 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
