magic
tech sky130A
magscale 1 2
timestamp 1672506959
<< metal2 >>
rect -4079 12180 -689 12502
rect -4079 11360 -3980 12180
rect -1520 11360 -689 12180
rect -4079 11002 -689 11360
tri -689 11002 811 12502 sw
tri -1311 9000 691 11002 ne
rect 691 10500 811 11002
tri 811 10500 1313 11002 sw
rect 691 10180 4024 10500
rect 691 9360 1480 10180
rect 3940 9360 4024 10180
rect 691 9000 4024 9360
rect 6408 400 15500 750
rect 6408 -440 6500 400
rect 7920 -440 15500 400
rect 6408 -750 15500 -440
tri -1311 -13004 691 -11002 se
rect 691 -11367 3925 -11002
rect 691 -12142 1392 -11367
rect 3841 -12142 3925 -11367
rect 691 -12502 3925 -12142
rect 691 -13004 811 -12502
tri 811 -13004 1313 -12502 nw
rect -4123 -13360 -689 -13004
rect -4123 -14135 -4031 -13360
rect -1582 -14135 -689 -13360
rect -4123 -14504 -689 -14135
tri -689 -14504 811 -13004 nw
<< via2 >>
rect -3980 11360 -1520 12180
rect 1480 9360 3940 10180
rect 6500 -440 7920 400
rect 1392 -12142 3841 -11367
rect -4031 -14135 -1582 -13360
<< metal3 >>
tri -7509 13004 -6009 14504 se
rect -6009 13004 6009 14504
tri 6009 13004 7509 14504 sw
tri -8642 11871 -7509 13004 se
rect -7509 12375 -6016 13004
tri -6016 12375 -5387 13004 nw
tri -5307 12375 -5180 12502 se
rect -5180 12375 -1739 12502
rect -7509 11871 -6725 12375
tri -9136 11377 -8642 11871 se
rect -8642 11666 -6725 11871
tri -6725 11666 -6016 12375 nw
tri -6016 11666 -5307 12375 se
rect -5307 12228 -1739 12375
tri -1739 12228 -1465 12502 sw
tri 562 12375 689 12502 se
rect 689 12375 5180 12502
tri 5180 12375 5307 12502 sw
tri 5387 12375 6016 13004 ne
rect 6016 12375 7509 13004
tri 415 12228 562 12375 se
rect 562 12255 5307 12375
tri 5307 12255 5427 12375 sw
tri 6016 12255 6136 12375 ne
rect 6136 12255 7509 12375
rect 562 12228 5427 12255
rect -5307 12180 -1453 12228
rect -5307 11666 -3980 12180
rect -8642 11377 -7302 11666
tri -10883 9630 -9136 11377 se
rect -9136 11089 -7302 11377
tri -7302 11089 -6725 11666 nw
tri -6305 11377 -6016 11666 se
rect -6016 11377 -3980 11666
tri -6593 11089 -6305 11377 se
rect -6305 11360 -3980 11377
rect -1520 11360 -1453 12180
rect -6305 11276 -1453 11360
rect -6305 11089 -1739 11276
rect -9136 10380 -8011 11089
tri -8011 10380 -7302 11089 nw
tri -7302 10380 -6593 11089 se
rect -6593 11002 -1739 11089
tri -1739 11002 -1465 11276 nw
rect -6593 10380 -5180 11002
tri -5180 10380 -4558 11002 nw
tri -1313 10500 415 12228 se
rect 415 11546 5427 12228
tri 5427 11546 6136 12255 sw
tri 6136 11546 6845 12255 ne
rect 6845 11546 7509 12255
tri 7509 11546 8967 13004 sw
rect 415 11002 6136 11546
rect 415 10500 433 11002
tri -4471 10380 -4351 10500 se
rect -4351 10380 433 10500
rect -9136 9868 -8523 10380
tri -8523 9868 -8011 10380 nw
tri -7814 9868 -7302 10380 se
rect -7302 9868 -5889 10380
rect -9136 9630 -9017 9868
tri -11139 9374 -10883 9630 se
rect -10883 9374 -9017 9630
tri -9017 9374 -8523 9868 nw
tri -8308 9374 -7814 9868 se
rect -7814 9671 -5889 9868
tri -5889 9671 -5180 10380 nw
tri -5180 9671 -4471 10380 se
rect -4471 10124 433 10380
tri 433 10124 1311 11002 nw
tri 4558 10500 5060 11002 ne
rect 5060 10837 6136 11002
tri 6136 10837 6845 11546 sw
tri 6845 10837 7554 11546 ne
rect 7554 10837 8967 11546
rect 5060 10500 6845 10837
tri 1410 10226 1684 10500 se
rect 1684 10253 4351 10500
tri 4351 10253 4598 10500 sw
tri 5060 10253 5307 10500 ne
rect 5307 10253 6845 10500
rect 1684 10226 4598 10253
rect 1410 10180 4598 10226
rect -4471 9671 -691 10124
rect -7814 9374 -6560 9671
tri -12382 8131 -11139 9374 se
rect -11139 8967 -9424 9374
tri -9424 8967 -9017 9374 nw
tri -8715 8967 -8308 9374 se
rect -8308 9000 -6560 9374
tri -6560 9000 -5889 9671 nw
tri -5851 9000 -5180 9671 se
rect -5180 9000 -691 9671
tri -691 9000 433 10124 nw
rect 1410 9360 1480 10180
rect 3940 9544 4598 10180
tri 4598 9544 5307 10253 sw
tri 5307 9544 6016 10253 ne
rect 6016 10133 6845 10253
tri 6845 10133 7549 10837 sw
tri 7554 10133 8258 10837 ne
rect 8258 10133 8967 10837
rect 6016 9544 7549 10133
rect 3940 9360 5307 9544
rect 1410 9274 5307 9360
tri 1410 9000 1684 9274 ne
rect 1684 9000 5307 9274
tri 5307 9000 5851 9544 sw
tri 6016 9000 6560 9544 ne
rect 6560 9424 7549 9544
tri 7549 9424 8258 10133 sw
tri 8258 9424 8967 10133 ne
tri 8967 9424 11089 11546 sw
rect 6560 9000 8258 9424
rect -8308 8967 -7182 9000
rect -11139 8258 -10133 8967
tri -10133 8258 -9424 8967 nw
tri -9424 8258 -8715 8967 se
rect -8715 8378 -7182 8967
tri -7182 8378 -6560 9000 nw
tri -6473 8378 -5851 9000 se
rect -5851 8378 -5427 9000
rect -8715 8258 -7429 8378
rect -11139 8131 -10260 8258
tri -10260 8131 -10133 8258 nw
tri -9551 8131 -9424 8258 se
rect -9424 8131 -7429 8258
tri -7429 8131 -7182 8378 nw
tri -6720 8131 -6473 8378 se
rect -6473 8131 -5427 8378
tri -14504 6009 -12382 8131 se
rect -12382 7422 -10969 8131
tri -10969 7422 -10260 8131 nw
tri -10260 7422 -9551 8131 se
rect -9551 7422 -8138 8131
tri -8138 7422 -7429 8131 nw
tri -7429 7422 -6720 8131 se
rect -6720 7422 -5427 8131
rect -12382 6845 -11546 7422
tri -11546 6845 -10969 7422 nw
tri -10837 6845 -10260 7422 se
rect -10260 6965 -8595 7422
tri -8595 6965 -8138 7422 nw
tri -7886 6965 -7429 7422 se
rect -7429 7302 -5427 7422
tri -5427 7302 -3729 9000 nw
tri 3729 7302 5427 9000 ne
rect 5427 8595 5851 9000
tri 5851 8595 6256 9000 sw
tri 6560 8595 6965 9000 ne
rect 6965 8715 8258 9000
tri 8258 8715 8967 9424 sw
tri 8967 8715 9676 9424 ne
rect 9676 8715 11089 9424
rect 6965 8595 8967 8715
rect 5427 8131 6256 8595
tri 6256 8131 6720 8595 sw
tri 6965 8131 7429 8595 ne
rect 7429 8131 8967 8595
rect 5427 7422 6720 8131
tri 6720 7422 7429 8131 sw
tri 7429 7422 8138 8131 ne
rect 8138 8011 8967 8131
tri 8967 8011 9671 8715 sw
tri 9676 8011 10380 8715 ne
rect 10380 8011 11089 8715
rect 8138 7422 9671 8011
rect 5427 7302 7429 7422
rect -7429 6965 -7342 7302
rect -10260 6845 -9304 6965
rect -12382 6136 -12255 6845
tri -12255 6136 -11546 6845 nw
tri -11546 6136 -10837 6845 se
rect -10837 6256 -9304 6845
tri -9304 6256 -8595 6965 nw
tri -8595 6256 -7886 6965 se
rect -7886 6256 -7342 6965
rect -10837 6136 -9551 6256
tri -12382 6009 -12255 6136 nw
rect -14504 -5889 -13004 6009
tri -13004 5387 -12382 6009 nw
tri -11793 5889 -11546 6136 se
rect -11546 6009 -9551 6136
tri -9551 6009 -9304 6256 nw
tri -8842 6009 -8595 6256 se
rect -8595 6009 -7342 6256
rect -11546 5889 -10173 6009
tri -12295 5387 -11793 5889 se
rect -11793 5387 -10173 5889
tri -10173 5387 -9551 6009 nw
tri -9464 5387 -8842 6009 se
rect -8842 5387 -7342 6009
tri -7342 5387 -5427 7302 nw
tri 5427 5387 7342 7302 ne
rect 7342 7182 7429 7302
tri 7429 7182 7669 7422 sw
tri 8138 7182 8378 7422 ne
rect 8378 7302 9671 7422
tri 9671 7302 10380 8011 sw
tri 10380 7302 11089 8011 ne
tri 11089 7302 13211 9424 sw
rect 8378 7182 10380 7302
rect 7342 6473 7669 7182
tri 7669 6473 8378 7182 sw
tri 8378 6473 9087 7182 ne
rect 9087 6593 10380 7182
tri 10380 6593 11089 7302 sw
tri 11089 6593 11798 7302 ne
rect 11798 6593 13211 7302
rect 9087 6473 11089 6593
rect 7342 6009 8378 6473
tri 8378 6009 8842 6473 sw
tri 9087 6009 9551 6473 ne
rect 9551 6009 11089 6473
rect 7342 5387 8842 6009
tri 8842 5387 9464 6009 sw
tri 9551 5387 10173 6009 ne
rect 10173 5889 11089 6009
tri 11089 5889 11793 6593 sw
tri 11798 5889 12502 6593 ne
rect 12502 6009 13211 6593
tri 13211 6009 14504 7302 sw
rect 12502 5889 14504 6009
rect 10173 5387 11793 5889
tri -12502 5180 -12295 5387 se
rect -12295 5180 -10500 5387
rect -12502 5060 -10500 5180
tri -10500 5060 -10173 5387 nw
tri -9791 5060 -9464 5387 se
rect -9464 5060 -9000 5387
rect -12502 -5060 -11002 5060
tri -11002 4558 -10500 5060 nw
tri -10500 4351 -9791 5060 se
rect -9791 4351 -9000 5060
rect -10500 750 -9000 4351
tri -9000 3729 -7342 5387 nw
tri 7342 3729 9000 5387 ne
rect 9000 5060 9464 5387
tri 9464 5060 9791 5387 sw
tri 10173 5060 10500 5387 ne
rect 10500 5180 11793 5387
tri 11793 5180 12502 5889 sw
tri 12502 5387 13004 5889 ne
rect 10500 5060 12502 5180
rect 9000 4351 9791 5060
tri 9791 4351 10500 5060 sw
tri 10500 4558 11002 5060 ne
rect -10500 400 8000 750
rect -10500 -440 6500 400
rect 7920 -440 8000 400
rect -10500 -750 8000 -440
rect -10500 -4351 -9000 -750
tri -11002 -5060 -10500 -4558 sw
tri -10500 -5060 -9791 -4351 ne
rect -9791 -5060 -9000 -4351
rect -12502 -5180 -10500 -5060
tri -13004 -5889 -12502 -5387 sw
tri -12502 -5889 -11793 -5180 ne
rect -11793 -5387 -10500 -5180
tri -10500 -5387 -10173 -5060 sw
tri -9791 -5387 -9464 -5060 ne
rect -9464 -5387 -9000 -5060
tri -9000 -5387 -7342 -3729 sw
tri 8171 -4558 9000 -3729 se
rect 9000 -4351 10500 4351
rect 9000 -4558 9791 -4351
rect -11793 -5889 -10173 -5387
rect -14504 -6009 -12502 -5889
tri -14504 -7302 -13211 -6009 ne
rect -13211 -6593 -12502 -6009
tri -12502 -6593 -11798 -5889 sw
tri -11793 -6593 -11089 -5889 ne
rect -11089 -6016 -10173 -5889
tri -10173 -6016 -9544 -5387 sw
tri -9464 -6016 -8835 -5387 ne
rect -8835 -6016 -7342 -5387
rect -11089 -6473 -9544 -6016
tri -9544 -6473 -9087 -6016 sw
tri -8835 -6473 -8378 -6016 ne
rect -8378 -6473 -7342 -6016
rect -11089 -6593 -9087 -6473
rect -13211 -7302 -11798 -6593
tri -11798 -7302 -11089 -6593 sw
tri -11089 -7302 -10380 -6593 ne
rect -10380 -7182 -9087 -6593
tri -9087 -7182 -8378 -6473 sw
tri -8378 -7182 -7669 -6473 ne
rect -7669 -7182 -7342 -6473
rect -10380 -7302 -8378 -7182
tri -13211 -9424 -11089 -7302 ne
tri -11089 -8011 -10380 -7302 sw
tri -10380 -8011 -9671 -7302 ne
rect -9671 -7422 -8378 -7302
tri -8378 -7422 -8138 -7182 sw
tri -7669 -7422 -7429 -7182 ne
rect -7429 -7302 -7342 -7182
tri -7342 -7302 -5427 -5387 sw
tri 6473 -6256 8171 -4558 se
rect 8171 -5060 9791 -4558
tri 9791 -5060 10500 -4351 nw
tri 10500 -5060 11002 -4558 se
rect 11002 -5060 12502 5060
rect 13004 3250 14504 5889
rect 13004 1750 15500 3250
rect 8171 -5387 9464 -5060
tri 9464 -5387 9791 -5060 nw
tri 10173 -5387 10500 -5060 se
rect 10500 -5180 12502 -5060
rect 10500 -5387 11793 -5180
rect 8171 -6016 8835 -5387
tri 8835 -6016 9464 -5387 nw
tri 9544 -6016 10173 -5387 se
rect 10173 -5889 11793 -5387
tri 11793 -5889 12502 -5180 nw
rect 13004 -3250 15500 -1750
tri 12502 -5889 13004 -5387 se
rect 13004 -5889 14504 -3250
rect 10173 -6016 11546 -5889
rect 8171 -6256 8595 -6016
tri 8595 -6256 8835 -6016 nw
tri 9304 -6256 9544 -6016 se
rect 9544 -6136 11546 -6016
tri 11546 -6136 11793 -5889 nw
tri 12255 -6136 12502 -5889 se
rect 12502 -6009 14504 -5889
rect 12502 -6136 14377 -6009
tri 14377 -6136 14504 -6009 nw
rect 9544 -6256 10837 -6136
tri 6256 -6473 6473 -6256 se
rect 6473 -6473 7886 -6256
tri 5427 -7302 6256 -6473 se
rect 6256 -6965 7886 -6473
tri 7886 -6965 8595 -6256 nw
tri 8595 -6965 9304 -6256 se
rect 9304 -6845 10837 -6256
tri 10837 -6845 11546 -6136 nw
tri 11546 -6845 12255 -6136 se
rect 9304 -6965 10253 -6845
rect 6256 -7302 7429 -6965
rect -7429 -7422 -5427 -7302
rect -9671 -8011 -8138 -7422
rect -11089 -8715 -10380 -8011
tri -10380 -8715 -9676 -8011 sw
tri -9671 -8715 -8967 -8011 ne
rect -8967 -8131 -8138 -8011
tri -8138 -8131 -7429 -7422 sw
tri -7429 -8131 -6720 -7422 ne
rect -6720 -8131 -5427 -7422
rect -8967 -8595 -7429 -8131
tri -7429 -8595 -6965 -8131 sw
tri -6720 -8595 -6256 -8131 ne
rect -6256 -8595 -5427 -8131
rect -8967 -8715 -6965 -8595
rect -11089 -9424 -9676 -8715
tri -9676 -9424 -8967 -8715 sw
tri -8967 -9424 -8258 -8715 ne
rect -8258 -9304 -6965 -8715
tri -6965 -9304 -6256 -8595 sw
tri -6256 -9304 -5547 -8595 ne
rect -5547 -9000 -5427 -8595
tri -5427 -9000 -3729 -7302 sw
tri 3729 -9000 5427 -7302 se
rect 5427 -7422 7429 -7302
tri 7429 -7422 7886 -6965 nw
tri 8138 -7422 8595 -6965 se
rect 8595 -7422 10253 -6965
rect 5427 -8131 6720 -7422
tri 6720 -8131 7429 -7422 nw
tri 7429 -8131 8138 -7422 se
rect 8138 -7429 10253 -7422
tri 10253 -7429 10837 -6845 nw
tri 10962 -7429 11546 -6845 se
rect 11546 -7429 12255 -6845
rect 8138 -8131 9544 -7429
rect 5427 -8378 6473 -8131
tri 6473 -8378 6720 -8131 nw
tri 7182 -8378 7429 -8131 se
rect 7429 -8138 9544 -8131
tri 9544 -8138 10253 -7429 nw
tri 10253 -8138 10962 -7429 se
rect 10962 -8138 12255 -7429
rect 7429 -8258 9424 -8138
tri 9424 -8258 9544 -8138 nw
tri 10133 -8258 10253 -8138 se
rect 10253 -8258 12255 -8138
tri 12255 -8258 14377 -6136 nw
rect 7429 -8378 8715 -8258
rect 5427 -9000 5764 -8378
rect -5547 -9087 5764 -9000
tri 5764 -9087 6473 -8378 nw
tri 6473 -9087 7182 -8378 se
rect 7182 -8967 8715 -8378
tri 8715 -8967 9424 -8258 nw
tri 9424 -8967 10133 -8258 se
rect 10133 -8967 10253 -8258
rect 7182 -9087 8131 -8967
rect -5547 -9304 5307 -9087
rect -8258 -9424 -6256 -9304
tri -11089 -11546 -8967 -9424 ne
tri -8967 -10133 -8258 -9424 sw
tri -8258 -10133 -7549 -9424 ne
rect -7549 -9544 -6256 -9424
tri -6256 -9544 -6016 -9304 sw
tri -5547 -9544 -5307 -9304 ne
rect -5307 -9544 5307 -9304
tri 5307 -9544 5764 -9087 nw
tri 6016 -9544 6473 -9087 se
rect 6473 -9544 8131 -9087
rect -7549 -10133 -6016 -9544
rect -8967 -10295 -8258 -10133
tri -8258 -10295 -8096 -10133 sw
tri -7549 -10295 -7387 -10133 ne
rect -7387 -10253 -6016 -10133
tri -6016 -10253 -5307 -9544 sw
tri -5307 -10253 -4598 -9544 ne
rect -4598 -10253 4598 -9544
tri 4598 -10253 5307 -9544 nw
tri 5307 -10253 6016 -9544 se
rect 6016 -9551 8131 -9544
tri 8131 -9551 8715 -8967 nw
tri 8840 -9551 9424 -8967 se
rect 9424 -9551 10253 -8967
rect 6016 -10253 7422 -9551
rect -7387 -10295 -5307 -10253
rect -8967 -11004 -8096 -10295
tri -8096 -11004 -7387 -10295 sw
tri -7387 -11004 -6678 -10295 ne
rect -6678 -10500 -5307 -10295
tri -5307 -10500 -5060 -10253 sw
tri -4598 -10500 -4351 -10253 ne
rect -4351 -10500 4351 -10253
tri 4351 -10500 4598 -10253 nw
tri 5060 -10500 5307 -10253 se
rect 5307 -10260 7422 -10253
tri 7422 -10260 8131 -9551 nw
tri 8131 -10260 8840 -9551 se
rect 8840 -10260 10253 -9551
tri 10253 -10260 12255 -8258 nw
rect 5307 -10380 7302 -10260
tri 7302 -10380 7422 -10260 nw
tri 8011 -10380 8131 -10260 se
rect 5307 -10500 6593 -10380
rect -6678 -11004 -5060 -10500
tri -5060 -11004 -4556 -10500 sw
tri 4558 -11002 5060 -10500 se
rect 5060 -11002 6593 -10500
rect -8967 -11546 -7387 -11004
tri -8967 -12502 -8011 -11546 ne
rect -8011 -11633 -7387 -11546
tri -7387 -11633 -6758 -11004 sw
tri -6678 -11633 -6049 -11004 ne
rect -6049 -11279 -689 -11004
tri -689 -11279 -414 -11004 sw
rect 1310 -11089 6593 -11002
tri 6593 -11089 7302 -10380 nw
tri 7302 -11089 8011 -10380 se
rect 8011 -11089 8131 -10380
rect 1310 -11279 6009 -11089
rect -6049 -11633 -414 -11279
rect -8011 -12255 -6758 -11633
tri -6758 -12255 -6136 -11633 sw
tri -6049 -12255 -5427 -11633 ne
rect -5427 -12255 -414 -11633
rect -8011 -12502 -6136 -12255
tri -6136 -12502 -5889 -12255 sw
tri -5427 -12502 -5180 -12255 ne
rect -5180 -12502 -414 -12255
tri -8011 -14504 -6009 -12502 ne
rect -6009 -13004 -5889 -12502
tri -5889 -13004 -5387 -12502 sw
tri -1313 -13004 -811 -12502 ne
rect -811 -13004 -414 -12502
tri -414 -13004 1311 -11279 sw
rect 1311 -11367 6009 -11279
rect 1311 -12142 1392 -11367
rect 3841 -11673 6009 -11367
tri 6009 -11673 6593 -11089 nw
tri 6718 -11673 7302 -11089 se
rect 7302 -11673 8131 -11089
rect 3841 -12142 5300 -11673
rect 1311 -12228 5300 -12142
tri 1311 -12502 1585 -12228 ne
rect 1585 -12382 5300 -12228
tri 5300 -12382 6009 -11673 nw
tri 6009 -12382 6718 -11673 se
rect 6718 -12382 8131 -11673
tri 8131 -12382 10253 -10260 nw
rect 1585 -12502 5180 -12382
tri 5180 -12502 5300 -12382 nw
tri 5387 -13004 6009 -12382 se
rect -6009 -13278 -1783 -13004
tri -1783 -13278 -1509 -13004 sw
rect -6009 -13360 -1509 -13278
rect -6009 -14135 -4031 -13360
rect -1582 -14135 -1509 -13360
rect -6009 -14230 -1509 -14135
rect -6009 -14504 -1783 -14230
tri -1783 -14504 -1509 -14230 nw
tri -811 -14504 689 -13004 ne
rect 689 -14504 6009 -13004
tri 6009 -14504 8131 -12382 nw
<< comment >>
tri -6009 6009 -2489 14504 ne
rect -2489 6009 2489 14504
tri 2489 6009 6009 14504 nw
tri -14504 2489 -6009 6009 sw
tri -2489 2489 -1031 6009 ne
rect -1031 2489 1031 6009
tri 1031 2490 2489 6009 nw
tri 6009 2490 14504 6009 se
rect -14504 427 -6009 2489
tri -6009 427 -1031 2489 sw
tri -1031 428 -177 2489 ne
rect -177 427 177 2489
tri 177 427 1031 2489 nw
tri 1031 427 6009 2489 se
rect 6009 427 14504 2490
rect -14504 73 -1031 427
tri -1031 73 -177 427 sw
tri -177 74 -31 427 ne
rect -31 73 30 427
tri 30 73 177 427 nw
tri 177 73 1031 427 se
rect 1031 73 14504 427
rect -14504 13 -177 73
tri -177 13 -31 73 sw
tri -31 13 -5 73 ne
rect -5 13 5 73
tri 5 13 30 73 nw
tri 30 13 177 73 se
rect 177 13 14504 73
rect -14504 2 -31 13
tri -31 2 -5 13 sw
tri -5 2 -1 13 ne
rect -1 2 1 13
tri 1 2 5 13 nw
tri 6 2 30 13 se
rect 30 2 14504 13
rect -14504 -2 -5 2
tri -5 0 -1 2 sw
tri -1 0 0 2 ne
tri 0 0 1 2 nw
tri 1 0 5 2 se
tri -5 -2 -1 0 nw
tri -1 -2 0 0 se
tri 0 -2 1 0 sw
tri 1 -2 5 0 ne
rect 5 -2 14504 2
rect -14504 -13 -30 -2
tri -30 -13 -5 -2 nw
tri -5 -13 -1 -2 se
rect -1 -12 1 -2
tri 1 -12 5 -2 sw
tri 5 -12 30 -2 ne
rect 30 -12 14504 -2
rect -1 -13 5 -12
rect -14504 -73 -177 -13
tri -177 -73 -30 -13 nw
tri -30 -73 -5 -13 se
rect -5 -73 5 -13
tri 5 -73 30 -12 sw
tri 30 -73 176 -12 ne
rect 176 -73 14504 -12
rect -14504 -427 -1031 -73
tri -1031 -427 -177 -73 nw
tri -177 -427 -30 -73 se
rect -30 -427 30 -73
tri 30 -427 177 -73 sw
tri 177 -427 1030 -73 ne
rect 1030 -427 14504 -73
rect -14504 -2489 -6009 -427
tri -6009 -2489 -1031 -427 nw
tri -1031 -2489 -177 -427 se
rect -177 -2489 177 -427
tri 177 -2489 1031 -427 sw
tri 1031 -2489 6008 -427 ne
rect 6008 -2489 14504 -427
tri -14504 -6009 -6009 -2489 nw
tri -2489 -6009 -1031 -2490 se
rect -1031 -6009 1031 -2489
tri 1031 -6009 2489 -2489 sw
tri 6009 -6009 14504 -2489 ne
tri -6009 -14504 -2489 -6009 se
rect -2489 -14504 2489 -6009
tri 2489 -14504 6009 -6009 sw
<< properties >>
string GDS_END 10489546
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_pr/gds/sky130_fd_pr.gds
string GDS_START 10482838
string gencell sky130_fd_pr__rf_test_coil1
string library sky130
string parameter m=1
string path 343.850 -150.225 343.850 -43.750 
<< end >>
