magic
tech sky130A
magscale 1 2
timestamp 1662478139
<< nwell >>
rect -246 -2281 246 2281
<< pmoslvt >>
rect -50 1862 50 2062
rect -50 1426 50 1626
rect -50 990 50 1190
rect -50 554 50 754
rect -50 118 50 318
rect -50 -318 50 -118
rect -50 -754 50 -554
rect -50 -1190 50 -990
rect -50 -1626 50 -1426
rect -50 -2062 50 -1862
<< pdiff >>
rect -108 2050 -50 2062
rect -108 1874 -96 2050
rect -62 1874 -50 2050
rect -108 1862 -50 1874
rect 50 2050 108 2062
rect 50 1874 62 2050
rect 96 1874 108 2050
rect 50 1862 108 1874
rect -108 1614 -50 1626
rect -108 1438 -96 1614
rect -62 1438 -50 1614
rect -108 1426 -50 1438
rect 50 1614 108 1626
rect 50 1438 62 1614
rect 96 1438 108 1614
rect 50 1426 108 1438
rect -108 1178 -50 1190
rect -108 1002 -96 1178
rect -62 1002 -50 1178
rect -108 990 -50 1002
rect 50 1178 108 1190
rect 50 1002 62 1178
rect 96 1002 108 1178
rect 50 990 108 1002
rect -108 742 -50 754
rect -108 566 -96 742
rect -62 566 -50 742
rect -108 554 -50 566
rect 50 742 108 754
rect 50 566 62 742
rect 96 566 108 742
rect 50 554 108 566
rect -108 306 -50 318
rect -108 130 -96 306
rect -62 130 -50 306
rect -108 118 -50 130
rect 50 306 108 318
rect 50 130 62 306
rect 96 130 108 306
rect 50 118 108 130
rect -108 -130 -50 -118
rect -108 -306 -96 -130
rect -62 -306 -50 -130
rect -108 -318 -50 -306
rect 50 -130 108 -118
rect 50 -306 62 -130
rect 96 -306 108 -130
rect 50 -318 108 -306
rect -108 -566 -50 -554
rect -108 -742 -96 -566
rect -62 -742 -50 -566
rect -108 -754 -50 -742
rect 50 -566 108 -554
rect 50 -742 62 -566
rect 96 -742 108 -566
rect 50 -754 108 -742
rect -108 -1002 -50 -990
rect -108 -1178 -96 -1002
rect -62 -1178 -50 -1002
rect -108 -1190 -50 -1178
rect 50 -1002 108 -990
rect 50 -1178 62 -1002
rect 96 -1178 108 -1002
rect 50 -1190 108 -1178
rect -108 -1438 -50 -1426
rect -108 -1614 -96 -1438
rect -62 -1614 -50 -1438
rect -108 -1626 -50 -1614
rect 50 -1438 108 -1426
rect 50 -1614 62 -1438
rect 96 -1614 108 -1438
rect 50 -1626 108 -1614
rect -108 -1874 -50 -1862
rect -108 -2050 -96 -1874
rect -62 -2050 -50 -1874
rect -108 -2062 -50 -2050
rect 50 -1874 108 -1862
rect 50 -2050 62 -1874
rect 96 -2050 108 -1874
rect 50 -2062 108 -2050
<< pdiffc >>
rect -96 1874 -62 2050
rect 62 1874 96 2050
rect -96 1438 -62 1614
rect 62 1438 96 1614
rect -96 1002 -62 1178
rect 62 1002 96 1178
rect -96 566 -62 742
rect 62 566 96 742
rect -96 130 -62 306
rect 62 130 96 306
rect -96 -306 -62 -130
rect 62 -306 96 -130
rect -96 -742 -62 -566
rect 62 -742 96 -566
rect -96 -1178 -62 -1002
rect 62 -1178 96 -1002
rect -96 -1614 -62 -1438
rect 62 -1614 96 -1438
rect -96 -2050 -62 -1874
rect 62 -2050 96 -1874
<< nsubdiff >>
rect -210 2211 -114 2245
rect 114 2211 210 2245
rect -210 2149 -176 2211
rect 176 2149 210 2211
rect -210 -2211 -176 -2149
rect 176 -2211 210 -2149
rect -210 -2245 -114 -2211
rect 114 -2245 210 -2211
<< nsubdiffcont >>
rect -114 2211 114 2245
rect -210 -2149 -176 2149
rect 176 -2149 210 2149
rect -114 -2245 114 -2211
<< poly >>
rect -50 2143 50 2159
rect -50 2109 -34 2143
rect 34 2109 50 2143
rect -50 2062 50 2109
rect -50 1815 50 1862
rect -50 1781 -34 1815
rect 34 1781 50 1815
rect -50 1765 50 1781
rect -50 1707 50 1723
rect -50 1673 -34 1707
rect 34 1673 50 1707
rect -50 1626 50 1673
rect -50 1379 50 1426
rect -50 1345 -34 1379
rect 34 1345 50 1379
rect -50 1329 50 1345
rect -50 1271 50 1287
rect -50 1237 -34 1271
rect 34 1237 50 1271
rect -50 1190 50 1237
rect -50 943 50 990
rect -50 909 -34 943
rect 34 909 50 943
rect -50 893 50 909
rect -50 835 50 851
rect -50 801 -34 835
rect 34 801 50 835
rect -50 754 50 801
rect -50 507 50 554
rect -50 473 -34 507
rect 34 473 50 507
rect -50 457 50 473
rect -50 399 50 415
rect -50 365 -34 399
rect 34 365 50 399
rect -50 318 50 365
rect -50 71 50 118
rect -50 37 -34 71
rect 34 37 50 71
rect -50 21 50 37
rect -50 -37 50 -21
rect -50 -71 -34 -37
rect 34 -71 50 -37
rect -50 -118 50 -71
rect -50 -365 50 -318
rect -50 -399 -34 -365
rect 34 -399 50 -365
rect -50 -415 50 -399
rect -50 -473 50 -457
rect -50 -507 -34 -473
rect 34 -507 50 -473
rect -50 -554 50 -507
rect -50 -801 50 -754
rect -50 -835 -34 -801
rect 34 -835 50 -801
rect -50 -851 50 -835
rect -50 -909 50 -893
rect -50 -943 -34 -909
rect 34 -943 50 -909
rect -50 -990 50 -943
rect -50 -1237 50 -1190
rect -50 -1271 -34 -1237
rect 34 -1271 50 -1237
rect -50 -1287 50 -1271
rect -50 -1345 50 -1329
rect -50 -1379 -34 -1345
rect 34 -1379 50 -1345
rect -50 -1426 50 -1379
rect -50 -1673 50 -1626
rect -50 -1707 -34 -1673
rect 34 -1707 50 -1673
rect -50 -1723 50 -1707
rect -50 -1781 50 -1765
rect -50 -1815 -34 -1781
rect 34 -1815 50 -1781
rect -50 -1862 50 -1815
rect -50 -2109 50 -2062
rect -50 -2143 -34 -2109
rect 34 -2143 50 -2109
rect -50 -2159 50 -2143
<< polycont >>
rect -34 2109 34 2143
rect -34 1781 34 1815
rect -34 1673 34 1707
rect -34 1345 34 1379
rect -34 1237 34 1271
rect -34 909 34 943
rect -34 801 34 835
rect -34 473 34 507
rect -34 365 34 399
rect -34 37 34 71
rect -34 -71 34 -37
rect -34 -399 34 -365
rect -34 -507 34 -473
rect -34 -835 34 -801
rect -34 -943 34 -909
rect -34 -1271 34 -1237
rect -34 -1379 34 -1345
rect -34 -1707 34 -1673
rect -34 -1815 34 -1781
rect -34 -2143 34 -2109
<< locali >>
rect -210 2211 -114 2245
rect 114 2211 210 2245
rect -210 2149 -176 2211
rect 176 2149 210 2211
rect -50 2109 -34 2143
rect 34 2109 50 2143
rect -96 2050 -62 2066
rect -96 1858 -62 1874
rect 62 2050 96 2066
rect 62 1858 96 1874
rect -50 1781 -34 1815
rect 34 1781 50 1815
rect -50 1673 -34 1707
rect 34 1673 50 1707
rect -96 1614 -62 1630
rect -96 1422 -62 1438
rect 62 1614 96 1630
rect 62 1422 96 1438
rect -50 1345 -34 1379
rect 34 1345 50 1379
rect -50 1237 -34 1271
rect 34 1237 50 1271
rect -96 1178 -62 1194
rect -96 986 -62 1002
rect 62 1178 96 1194
rect 62 986 96 1002
rect -50 909 -34 943
rect 34 909 50 943
rect -50 801 -34 835
rect 34 801 50 835
rect -96 742 -62 758
rect -96 550 -62 566
rect 62 742 96 758
rect 62 550 96 566
rect -50 473 -34 507
rect 34 473 50 507
rect -50 365 -34 399
rect 34 365 50 399
rect -96 306 -62 322
rect -96 114 -62 130
rect 62 306 96 322
rect 62 114 96 130
rect -50 37 -34 71
rect 34 37 50 71
rect -50 -71 -34 -37
rect 34 -71 50 -37
rect -96 -130 -62 -114
rect -96 -322 -62 -306
rect 62 -130 96 -114
rect 62 -322 96 -306
rect -50 -399 -34 -365
rect 34 -399 50 -365
rect -50 -507 -34 -473
rect 34 -507 50 -473
rect -96 -566 -62 -550
rect -96 -758 -62 -742
rect 62 -566 96 -550
rect 62 -758 96 -742
rect -50 -835 -34 -801
rect 34 -835 50 -801
rect -50 -943 -34 -909
rect 34 -943 50 -909
rect -96 -1002 -62 -986
rect -96 -1194 -62 -1178
rect 62 -1002 96 -986
rect 62 -1194 96 -1178
rect -50 -1271 -34 -1237
rect 34 -1271 50 -1237
rect -50 -1379 -34 -1345
rect 34 -1379 50 -1345
rect -96 -1438 -62 -1422
rect -96 -1630 -62 -1614
rect 62 -1438 96 -1422
rect 62 -1630 96 -1614
rect -50 -1707 -34 -1673
rect 34 -1707 50 -1673
rect -50 -1815 -34 -1781
rect 34 -1815 50 -1781
rect -96 -1874 -62 -1858
rect -96 -2066 -62 -2050
rect 62 -1874 96 -1858
rect 62 -2066 96 -2050
rect -50 -2143 -34 -2109
rect 34 -2143 50 -2109
rect -210 -2211 -176 -2149
rect 176 -2211 210 -2149
rect -210 -2245 -114 -2211
rect 114 -2245 210 -2211
<< viali >>
rect -34 2109 34 2143
rect -96 1874 -62 2050
rect 62 1874 96 2050
rect -34 1781 34 1815
rect -34 1673 34 1707
rect -96 1438 -62 1614
rect 62 1438 96 1614
rect -34 1345 34 1379
rect -34 1237 34 1271
rect -96 1002 -62 1178
rect 62 1002 96 1178
rect -34 909 34 943
rect -34 801 34 835
rect -96 566 -62 742
rect 62 566 96 742
rect -34 473 34 507
rect -34 365 34 399
rect -96 130 -62 306
rect 62 130 96 306
rect -34 37 34 71
rect -34 -71 34 -37
rect -96 -306 -62 -130
rect 62 -306 96 -130
rect -34 -399 34 -365
rect -34 -507 34 -473
rect -96 -742 -62 -566
rect 62 -742 96 -566
rect -34 -835 34 -801
rect -34 -943 34 -909
rect -96 -1178 -62 -1002
rect 62 -1178 96 -1002
rect -34 -1271 34 -1237
rect -34 -1379 34 -1345
rect -96 -1614 -62 -1438
rect 62 -1614 96 -1438
rect -34 -1707 34 -1673
rect -34 -1815 34 -1781
rect -96 -2050 -62 -1874
rect 62 -2050 96 -1874
rect -34 -2143 34 -2109
<< metal1 >>
rect -46 2143 46 2149
rect -46 2109 -34 2143
rect 34 2109 46 2143
rect -46 2103 46 2109
rect -102 2050 -56 2062
rect -102 1874 -96 2050
rect -62 1874 -56 2050
rect -102 1862 -56 1874
rect 56 2050 102 2062
rect 56 1874 62 2050
rect 96 1874 102 2050
rect 56 1862 102 1874
rect -46 1815 46 1821
rect -46 1781 -34 1815
rect 34 1781 46 1815
rect -46 1775 46 1781
rect -46 1707 46 1713
rect -46 1673 -34 1707
rect 34 1673 46 1707
rect -46 1667 46 1673
rect -102 1614 -56 1626
rect -102 1438 -96 1614
rect -62 1438 -56 1614
rect -102 1426 -56 1438
rect 56 1614 102 1626
rect 56 1438 62 1614
rect 96 1438 102 1614
rect 56 1426 102 1438
rect -46 1379 46 1385
rect -46 1345 -34 1379
rect 34 1345 46 1379
rect -46 1339 46 1345
rect -46 1271 46 1277
rect -46 1237 -34 1271
rect 34 1237 46 1271
rect -46 1231 46 1237
rect -102 1178 -56 1190
rect -102 1002 -96 1178
rect -62 1002 -56 1178
rect -102 990 -56 1002
rect 56 1178 102 1190
rect 56 1002 62 1178
rect 96 1002 102 1178
rect 56 990 102 1002
rect -46 943 46 949
rect -46 909 -34 943
rect 34 909 46 943
rect -46 903 46 909
rect -46 835 46 841
rect -46 801 -34 835
rect 34 801 46 835
rect -46 795 46 801
rect -102 742 -56 754
rect -102 566 -96 742
rect -62 566 -56 742
rect -102 554 -56 566
rect 56 742 102 754
rect 56 566 62 742
rect 96 566 102 742
rect 56 554 102 566
rect -46 507 46 513
rect -46 473 -34 507
rect 34 473 46 507
rect -46 467 46 473
rect -46 399 46 405
rect -46 365 -34 399
rect 34 365 46 399
rect -46 359 46 365
rect -102 306 -56 318
rect -102 130 -96 306
rect -62 130 -56 306
rect -102 118 -56 130
rect 56 306 102 318
rect 56 130 62 306
rect 96 130 102 306
rect 56 118 102 130
rect -46 71 46 77
rect -46 37 -34 71
rect 34 37 46 71
rect -46 31 46 37
rect -46 -37 46 -31
rect -46 -71 -34 -37
rect 34 -71 46 -37
rect -46 -77 46 -71
rect -102 -130 -56 -118
rect -102 -306 -96 -130
rect -62 -306 -56 -130
rect -102 -318 -56 -306
rect 56 -130 102 -118
rect 56 -306 62 -130
rect 96 -306 102 -130
rect 56 -318 102 -306
rect -46 -365 46 -359
rect -46 -399 -34 -365
rect 34 -399 46 -365
rect -46 -405 46 -399
rect -46 -473 46 -467
rect -46 -507 -34 -473
rect 34 -507 46 -473
rect -46 -513 46 -507
rect -102 -566 -56 -554
rect -102 -742 -96 -566
rect -62 -742 -56 -566
rect -102 -754 -56 -742
rect 56 -566 102 -554
rect 56 -742 62 -566
rect 96 -742 102 -566
rect 56 -754 102 -742
rect -46 -801 46 -795
rect -46 -835 -34 -801
rect 34 -835 46 -801
rect -46 -841 46 -835
rect -46 -909 46 -903
rect -46 -943 -34 -909
rect 34 -943 46 -909
rect -46 -949 46 -943
rect -102 -1002 -56 -990
rect -102 -1178 -96 -1002
rect -62 -1178 -56 -1002
rect -102 -1190 -56 -1178
rect 56 -1002 102 -990
rect 56 -1178 62 -1002
rect 96 -1178 102 -1002
rect 56 -1190 102 -1178
rect -46 -1237 46 -1231
rect -46 -1271 -34 -1237
rect 34 -1271 46 -1237
rect -46 -1277 46 -1271
rect -46 -1345 46 -1339
rect -46 -1379 -34 -1345
rect 34 -1379 46 -1345
rect -46 -1385 46 -1379
rect -102 -1438 -56 -1426
rect -102 -1614 -96 -1438
rect -62 -1614 -56 -1438
rect -102 -1626 -56 -1614
rect 56 -1438 102 -1426
rect 56 -1614 62 -1438
rect 96 -1614 102 -1438
rect 56 -1626 102 -1614
rect -46 -1673 46 -1667
rect -46 -1707 -34 -1673
rect 34 -1707 46 -1673
rect -46 -1713 46 -1707
rect -46 -1781 46 -1775
rect -46 -1815 -34 -1781
rect 34 -1815 46 -1781
rect -46 -1821 46 -1815
rect -102 -1874 -56 -1862
rect -102 -2050 -96 -1874
rect -62 -2050 -56 -1874
rect -102 -2062 -56 -2050
rect 56 -1874 102 -1862
rect 56 -2050 62 -1874
rect 96 -2050 102 -1874
rect 56 -2062 102 -2050
rect -46 -2109 46 -2103
rect -46 -2143 -34 -2109
rect 34 -2143 46 -2109
rect -46 -2149 46 -2143
<< properties >>
string FIXED_BBOX -193 -2228 193 2228
string gencell sky130_fd_pr__pfet_01v8_lvt
string library sky130
string parameters w 1.0 l 0.5 m 10 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.35 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
