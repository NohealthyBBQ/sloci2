magic
tech sky130A
magscale 1 2
timestamp 1672460674
<< locali >>
rect -14000 -57650 -13940 -57640
rect -14000 -57690 -13990 -57650
rect -13950 -57690 -13940 -57650
rect -14000 -57700 -13940 -57690
<< viali >>
rect -13990 -57690 -13950 -57650
<< metal1 >>
rect -14303 -57650 -13881 -57599
rect -14303 -57690 -13990 -57650
rect -13950 -57690 -13881 -57650
rect -14303 -57950 -13881 -57690
rect -14303 -58050 -14250 -57950
rect -14150 -58050 -13881 -57950
rect -14303 -58103 -13881 -58050
<< via1 >>
rect -14250 -58050 -14150 -57950
<< metal2 >>
rect -14303 -57950 -13881 -57599
rect -14303 -58050 -14250 -57950
rect -14150 -58050 -13881 -57950
rect -14303 -58103 -13881 -58050
<< via2 >>
rect -14250 -58050 -14150 -57950
<< metal3 >>
rect -17920 -57950 19840 35200
rect -17920 -58050 -14250 -57950
rect -14150 -58050 19840 -57950
rect -17920 -62080 19840 -58050
<< metal4 >>
rect 960 17560 1280 17600
rect 960 17320 1000 17560
rect 1240 17320 1280 17560
rect 960 -13160 1280 17320
rect 960 -13400 1000 -13160
rect 1240 -13400 1280 -13160
rect 960 -37480 1280 -13400
rect 960 -37720 1000 -37480
rect 1240 -37720 1280 -37480
rect 960 -52520 1280 -37720
rect 960 -52760 1000 -52520
rect 1240 -52760 1280 -52520
rect 960 -52800 1280 -52760
<< via4 >>
rect 1000 17320 1240 17560
rect 1000 -13400 1240 -13160
rect 1000 -37720 1240 -37480
rect 1000 -52760 1240 -52520
<< metal5 >>
rect -8640 26880 10560 27200
rect -8640 8000 -8320 26880
rect -8000 26240 9920 26560
rect -8000 8640 -7680 26240
rect -7360 25600 9280 25920
rect -7360 9280 -7040 25600
rect -6720 24960 8640 25280
rect -6720 9920 -6400 24960
rect -6080 24320 8000 24640
rect -6080 10560 -5760 24320
rect -5440 23680 7360 24000
rect -5440 11200 -5120 23680
rect -4800 23040 6720 23360
rect -4800 11840 -4480 23040
rect -4160 22400 6080 22720
rect -4160 12480 -3840 22400
rect -3520 21760 5440 22080
rect -3520 13120 -3200 21760
rect -2880 21120 4800 21440
rect -2880 13760 -2560 21120
rect -2240 20480 4160 20800
rect -2240 14400 -1920 20480
rect -1600 19840 3520 20160
rect -1600 15040 -1280 19840
rect -960 19200 2880 19520
rect -960 15680 -640 19200
rect -320 18560 2240 18880
rect -320 16320 0 18560
rect 320 17920 1600 18240
rect 320 16960 640 17920
rect 1280 17600 1600 17920
rect 960 17560 1600 17600
rect 960 17320 1000 17560
rect 1240 17320 1600 17560
rect 960 17280 1600 17320
rect 1920 16960 2240 18560
rect 320 16640 2240 16960
rect 2560 16320 2880 19200
rect -320 16000 2880 16320
rect 3200 15680 3520 19840
rect -960 15360 3520 15680
rect 3840 15040 4160 20480
rect -1600 14720 4160 15040
rect 4480 14400 4800 21120
rect -2240 14080 4800 14400
rect 5120 13760 5440 21760
rect -2880 13440 5440 13760
rect 5760 13120 6080 22400
rect -3520 12800 6080 13120
rect 6400 12480 6720 23040
rect -4160 12160 6720 12480
rect 7040 11840 7360 23680
rect -4800 11520 7360 11840
rect 7680 11200 8000 24320
rect -5440 10880 8000 11200
rect 8320 10560 8640 24960
rect -6080 10240 8640 10560
rect 8960 9920 9280 25600
rect -6720 9600 9280 9920
rect 9600 9280 9920 26240
rect -7360 8960 9920 9280
rect 10240 8640 10560 26880
rect -8000 8320 10560 8640
rect -8640 7680 10880 8000
rect -6720 -5760 8640 -5440
rect -6720 -20800 -6400 -5760
rect -6080 -6400 8000 -6080
rect -6080 -20160 -5760 -6400
rect -5440 -7040 7360 -6720
rect -5440 -19520 -5120 -7040
rect -4800 -7680 6720 -7360
rect -4800 -18880 -4480 -7680
rect -4160 -8320 6080 -8000
rect -4160 -18240 -3840 -8320
rect -3520 -8960 5440 -8640
rect -3520 -17600 -3200 -8960
rect -2880 -9600 4800 -9280
rect -2880 -16960 -2560 -9600
rect -2240 -10240 4160 -9920
rect -2240 -16320 -1920 -10240
rect -1600 -10880 3520 -10560
rect -1600 -15680 -1280 -10880
rect -960 -11520 2880 -11200
rect -960 -15040 -640 -11520
rect -320 -12160 2240 -11840
rect -320 -14400 0 -12160
rect 320 -12800 1600 -12480
rect 320 -13760 640 -12800
rect 1280 -13120 1600 -12800
rect 960 -13160 1600 -13120
rect 960 -13400 1000 -13160
rect 1240 -13400 1600 -13160
rect 960 -13440 1600 -13400
rect 1920 -13760 2240 -12160
rect 320 -14080 2240 -13760
rect 2560 -14400 2880 -11520
rect -320 -14720 2880 -14400
rect 3200 -15040 3520 -10880
rect -960 -15360 3520 -15040
rect 3840 -15680 4160 -10240
rect -1600 -16000 4160 -15680
rect 4480 -16320 4800 -9600
rect -2240 -16640 4800 -16320
rect 5120 -16960 5440 -8960
rect -2880 -17280 5440 -16960
rect 5760 -17600 6080 -8320
rect -3520 -17920 6080 -17600
rect 6400 -18240 6720 -7680
rect -4160 -18560 6720 -18240
rect 7040 -18880 7360 -7040
rect -4800 -19200 7360 -18880
rect 7680 -19520 8000 -6400
rect -5440 -19840 8000 -19520
rect 8320 -20160 8640 -5760
rect -6080 -20480 8640 -20160
rect -6720 -21120 8960 -20800
rect -4160 -32640 6080 -32320
rect -4160 -42560 -3840 -32640
rect -3520 -33280 5440 -32960
rect -3520 -41920 -3200 -33280
rect -2880 -33920 4800 -33600
rect -2880 -41280 -2560 -33920
rect -2240 -34560 4160 -34240
rect -2240 -40640 -1920 -34560
rect -1600 -35200 3520 -34880
rect -1600 -40000 -1280 -35200
rect -960 -35840 2880 -35520
rect -960 -39360 -640 -35840
rect -320 -36480 2240 -36160
rect -320 -38720 0 -36480
rect 320 -37120 1600 -36800
rect 320 -38080 640 -37120
rect 1280 -37440 1600 -37120
rect 960 -37480 1600 -37440
rect 960 -37720 1000 -37480
rect 1240 -37720 1600 -37480
rect 960 -37760 1600 -37720
rect 1920 -38080 2240 -36480
rect 320 -38400 2240 -38080
rect 2560 -38720 2880 -35840
rect -320 -39040 2880 -38720
rect 3200 -39360 3520 -35200
rect -960 -39680 3520 -39360
rect 3840 -40000 4160 -34560
rect -1600 -40320 4160 -40000
rect 4480 -40640 4800 -33920
rect -2240 -40960 4800 -40640
rect 5120 -41280 5440 -33280
rect -2880 -41600 5440 -41280
rect 5760 -41920 6080 -32640
rect -3520 -42240 6080 -41920
rect -4160 -42880 6400 -42560
rect -1600 -50240 3520 -49920
rect -1600 -55040 -1280 -50240
rect -960 -50880 2880 -50560
rect -960 -54400 -640 -50880
rect -320 -51520 2240 -51200
rect -320 -53760 0 -51520
rect 320 -52160 1600 -51840
rect 320 -53120 640 -52160
rect 1280 -52480 1600 -52160
rect 960 -52520 1600 -52480
rect 960 -52760 1000 -52520
rect 1240 -52760 1600 -52520
rect 960 -52800 1600 -52760
rect 1920 -53120 2240 -51520
rect 320 -53440 2240 -53120
rect 2560 -53760 2880 -50880
rect -320 -54080 2880 -53760
rect 3200 -54400 3520 -50240
rect -960 -54720 3520 -54400
rect -1600 -55360 3840 -55040
use sky130_fd_pr__nfet_01v8_EDB9KC  sky130_fd_pr__nfet_01v8_EDB9KC_0
timestamp 1672460213
transform 1 0 -14092 0 1 -57851
box -211 -252 211 252
<< end >>
