magic
tech sky130A
magscale 1 2
timestamp 1662690363
<< error_p >>
rect -159 181 -97 187
rect -31 181 31 187
rect 97 181 159 187
rect -159 147 -147 181
rect -31 147 -19 181
rect 97 147 109 181
rect -159 141 -97 147
rect -31 141 31 147
rect 97 141 159 147
rect -159 -147 -97 -141
rect -31 -147 31 -141
rect 97 -147 159 -141
rect -159 -181 -147 -147
rect -31 -181 -19 -147
rect 97 -181 109 -147
rect -159 -187 -97 -181
rect -31 -187 31 -181
rect 97 -187 159 -181
<< nwell >>
rect -359 -319 359 319
<< pmoslvt >>
rect -163 -100 -93 100
rect -35 -100 35 100
rect 93 -100 163 100
<< pdiff >>
rect -221 88 -163 100
rect -221 -88 -209 88
rect -175 -88 -163 88
rect -221 -100 -163 -88
rect -93 88 -35 100
rect -93 -88 -81 88
rect -47 -88 -35 88
rect -93 -100 -35 -88
rect 35 88 93 100
rect 35 -88 47 88
rect 81 -88 93 88
rect 35 -100 93 -88
rect 163 88 221 100
rect 163 -88 175 88
rect 209 -88 221 88
rect 163 -100 221 -88
<< pdiffc >>
rect -209 -88 -175 88
rect -81 -88 -47 88
rect 47 -88 81 88
rect 175 -88 209 88
<< nsubdiff >>
rect -323 249 -227 283
rect 227 249 323 283
rect -323 187 -289 249
rect 289 187 323 249
rect -323 -249 -289 -187
rect 289 -249 323 -187
rect -323 -283 -227 -249
rect 227 -283 323 -249
<< nsubdiffcont >>
rect -227 249 227 283
rect -323 -187 -289 187
rect 289 -187 323 187
rect -227 -283 227 -249
<< poly >>
rect -163 181 -93 197
rect -163 147 -147 181
rect -109 147 -93 181
rect -163 100 -93 147
rect -35 181 35 197
rect -35 147 -19 181
rect 19 147 35 181
rect -35 100 35 147
rect 93 181 163 197
rect 93 147 109 181
rect 147 147 163 181
rect 93 100 163 147
rect -163 -147 -93 -100
rect -163 -181 -147 -147
rect -109 -181 -93 -147
rect -163 -197 -93 -181
rect -35 -147 35 -100
rect -35 -181 -19 -147
rect 19 -181 35 -147
rect -35 -197 35 -181
rect 93 -147 163 -100
rect 93 -181 109 -147
rect 147 -181 163 -147
rect 93 -197 163 -181
<< polycont >>
rect -147 147 -109 181
rect -19 147 19 181
rect 109 147 147 181
rect -147 -181 -109 -147
rect -19 -181 19 -147
rect 109 -181 147 -147
<< locali >>
rect -323 249 -227 283
rect 227 249 323 283
rect -323 187 -289 249
rect 289 187 323 249
rect -163 147 -147 181
rect -109 147 -93 181
rect -35 147 -19 181
rect 19 147 35 181
rect 93 147 109 181
rect 147 147 163 181
rect -209 88 -175 104
rect -209 -104 -175 -88
rect -81 88 -47 104
rect -81 -104 -47 -88
rect 47 88 81 104
rect 47 -104 81 -88
rect 175 88 209 104
rect 175 -104 209 -88
rect -163 -181 -147 -147
rect -109 -181 -93 -147
rect -35 -181 -19 -147
rect 19 -181 35 -147
rect 93 -181 109 -147
rect 147 -181 163 -147
rect -323 -249 -289 -187
rect 289 -249 323 -187
rect -323 -283 -227 -249
rect 227 -283 323 -249
<< viali >>
rect -147 147 -109 181
rect -19 147 19 181
rect 109 147 147 181
rect -209 -88 -175 88
rect -81 -88 -47 88
rect 47 -88 81 88
rect 175 -88 209 88
rect -147 -181 -109 -147
rect -19 -181 19 -147
rect 109 -181 147 -147
<< metal1 >>
rect -159 181 -97 187
rect -159 147 -147 181
rect -109 147 -97 181
rect -159 141 -97 147
rect -31 181 31 187
rect -31 147 -19 181
rect 19 147 31 181
rect -31 141 31 147
rect 97 181 159 187
rect 97 147 109 181
rect 147 147 159 181
rect 97 141 159 147
rect -215 88 -169 100
rect -215 -88 -209 88
rect -175 -88 -169 88
rect -215 -100 -169 -88
rect -87 88 -41 100
rect -87 -88 -81 88
rect -47 -88 -41 88
rect -87 -100 -41 -88
rect 41 88 87 100
rect 41 -88 47 88
rect 81 -88 87 88
rect 41 -100 87 -88
rect 169 88 215 100
rect 169 -88 175 88
rect 209 -88 215 88
rect 169 -100 215 -88
rect -159 -147 -97 -141
rect -159 -181 -147 -147
rect -109 -181 -97 -147
rect -159 -187 -97 -181
rect -31 -147 31 -141
rect -31 -181 -19 -147
rect 19 -181 31 -147
rect -31 -187 31 -181
rect 97 -147 159 -141
rect 97 -181 109 -147
rect 147 -181 159 -147
rect 97 -187 159 -181
<< properties >>
string FIXED_BBOX -306 -266 306 266
string gencell sky130_fd_pr__pfet_01v8_lvt
string library sky130
string parameters w 1 l 0.35 m 1 nf 3 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.35 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
