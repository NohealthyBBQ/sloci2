** sch_path: /home/zexi/sloci/design/misc/single_mos_lvs/nfet_nf1_m8.sch
**.subckt nfet_nf1_m8 G S B D
*.ipin G
*.iopin S
*.iopin B
*.opin D
XM1 D G S B sky130_fd_pr__nfet_01v8_lvt L=1 W=2 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=8 m=8
**.ends
.end
