magic
tech sky130A
timestamp 1671767400
<< pwell >>
rect -1524 -155 1523 155
<< nmoslvt >>
rect -1424 -50 -1409 50
rect -1376 -50 -1361 50
rect -1328 -50 -1313 50
rect -1280 -50 -1265 50
rect -1232 -50 -1217 50
rect -1184 -50 -1169 50
rect -1136 -50 -1121 50
rect -1088 -50 -1073 50
rect -1040 -50 -1025 50
rect -992 -50 -977 50
rect -944 -50 -929 50
rect -896 -50 -881 50
rect -848 -50 -833 50
rect -800 -50 -785 50
rect -752 -50 -737 50
rect -704 -50 -689 50
rect -656 -50 -641 50
rect -608 -50 -593 50
rect -560 -50 -545 50
rect -512 -50 -497 50
rect -464 -50 -449 50
rect -416 -50 -401 50
rect -368 -50 -353 50
rect -320 -50 -305 50
rect -272 -50 -257 50
rect -224 -50 -209 50
rect -176 -50 -161 50
rect -128 -50 -113 50
rect -80 -50 -65 50
rect -32 -50 -17 50
rect 16 -50 31 50
rect 64 -50 79 50
rect 112 -50 127 50
rect 160 -50 175 50
rect 208 -50 223 50
rect 256 -50 271 50
rect 304 -50 319 50
rect 352 -50 367 50
rect 400 -50 415 50
rect 448 -50 463 50
rect 496 -50 511 50
rect 544 -50 559 50
rect 592 -50 607 50
rect 640 -50 655 50
rect 688 -50 703 50
rect 736 -50 751 50
rect 784 -50 799 50
rect 832 -50 847 50
rect 880 -50 895 50
rect 928 -50 943 50
rect 976 -50 991 50
rect 1024 -50 1039 50
rect 1072 -50 1087 50
rect 1120 -50 1135 50
rect 1168 -50 1183 50
rect 1216 -50 1231 50
rect 1264 -50 1279 50
rect 1312 -50 1327 50
rect 1360 -50 1375 50
rect 1408 -50 1423 50
<< ndiff >>
rect -1455 44 -1424 50
rect -1455 -44 -1449 44
rect -1432 -44 -1424 44
rect -1455 -50 -1424 -44
rect -1409 44 -1376 50
rect -1409 -44 -1401 44
rect -1384 -44 -1376 44
rect -1409 -50 -1376 -44
rect -1361 44 -1328 50
rect -1361 -44 -1353 44
rect -1336 -44 -1328 44
rect -1361 -50 -1328 -44
rect -1313 44 -1280 50
rect -1313 -44 -1305 44
rect -1288 -44 -1280 44
rect -1313 -50 -1280 -44
rect -1265 44 -1232 50
rect -1265 -44 -1257 44
rect -1240 -44 -1232 44
rect -1265 -50 -1232 -44
rect -1217 44 -1184 50
rect -1217 -44 -1209 44
rect -1192 -44 -1184 44
rect -1217 -50 -1184 -44
rect -1169 44 -1136 50
rect -1169 -44 -1161 44
rect -1144 -44 -1136 44
rect -1169 -50 -1136 -44
rect -1121 44 -1088 50
rect -1121 -44 -1113 44
rect -1096 -44 -1088 44
rect -1121 -50 -1088 -44
rect -1073 44 -1040 50
rect -1073 -44 -1065 44
rect -1048 -44 -1040 44
rect -1073 -50 -1040 -44
rect -1025 44 -992 50
rect -1025 -44 -1017 44
rect -1000 -44 -992 44
rect -1025 -50 -992 -44
rect -977 44 -944 50
rect -977 -44 -969 44
rect -952 -44 -944 44
rect -977 -50 -944 -44
rect -929 44 -896 50
rect -929 -44 -921 44
rect -904 -44 -896 44
rect -929 -50 -896 -44
rect -881 44 -848 50
rect -881 -44 -873 44
rect -856 -44 -848 44
rect -881 -50 -848 -44
rect -833 44 -800 50
rect -833 -44 -825 44
rect -808 -44 -800 44
rect -833 -50 -800 -44
rect -785 44 -752 50
rect -785 -44 -777 44
rect -760 -44 -752 44
rect -785 -50 -752 -44
rect -737 44 -704 50
rect -737 -44 -729 44
rect -712 -44 -704 44
rect -737 -50 -704 -44
rect -689 44 -656 50
rect -689 -44 -681 44
rect -664 -44 -656 44
rect -689 -50 -656 -44
rect -641 44 -608 50
rect -641 -44 -633 44
rect -616 -44 -608 44
rect -641 -50 -608 -44
rect -593 44 -560 50
rect -593 -44 -585 44
rect -568 -44 -560 44
rect -593 -50 -560 -44
rect -545 44 -512 50
rect -545 -44 -537 44
rect -520 -44 -512 44
rect -545 -50 -512 -44
rect -497 44 -464 50
rect -497 -44 -489 44
rect -472 -44 -464 44
rect -497 -50 -464 -44
rect -449 44 -416 50
rect -449 -44 -441 44
rect -424 -44 -416 44
rect -449 -50 -416 -44
rect -401 44 -368 50
rect -401 -44 -393 44
rect -376 -44 -368 44
rect -401 -50 -368 -44
rect -353 44 -320 50
rect -353 -44 -345 44
rect -328 -44 -320 44
rect -353 -50 -320 -44
rect -305 44 -272 50
rect -305 -44 -297 44
rect -280 -44 -272 44
rect -305 -50 -272 -44
rect -257 44 -224 50
rect -257 -44 -249 44
rect -232 -44 -224 44
rect -257 -50 -224 -44
rect -209 44 -176 50
rect -209 -44 -201 44
rect -184 -44 -176 44
rect -209 -50 -176 -44
rect -161 44 -128 50
rect -161 -44 -153 44
rect -136 -44 -128 44
rect -161 -50 -128 -44
rect -113 44 -80 50
rect -113 -44 -105 44
rect -88 -44 -80 44
rect -113 -50 -80 -44
rect -65 44 -32 50
rect -65 -44 -57 44
rect -40 -44 -32 44
rect -65 -50 -32 -44
rect -17 44 16 50
rect -17 -44 -9 44
rect 8 -44 16 44
rect -17 -50 16 -44
rect 31 44 64 50
rect 31 -44 39 44
rect 56 -44 64 44
rect 31 -50 64 -44
rect 79 44 112 50
rect 79 -44 87 44
rect 104 -44 112 44
rect 79 -50 112 -44
rect 127 44 160 50
rect 127 -44 135 44
rect 152 -44 160 44
rect 127 -50 160 -44
rect 175 44 208 50
rect 175 -44 183 44
rect 200 -44 208 44
rect 175 -50 208 -44
rect 223 44 256 50
rect 223 -44 231 44
rect 248 -44 256 44
rect 223 -50 256 -44
rect 271 44 304 50
rect 271 -44 279 44
rect 296 -44 304 44
rect 271 -50 304 -44
rect 319 44 352 50
rect 319 -44 327 44
rect 344 -44 352 44
rect 319 -50 352 -44
rect 367 44 400 50
rect 367 -44 375 44
rect 392 -44 400 44
rect 367 -50 400 -44
rect 415 44 448 50
rect 415 -44 423 44
rect 440 -44 448 44
rect 415 -50 448 -44
rect 463 44 496 50
rect 463 -44 471 44
rect 488 -44 496 44
rect 463 -50 496 -44
rect 511 44 544 50
rect 511 -44 519 44
rect 536 -44 544 44
rect 511 -50 544 -44
rect 559 44 592 50
rect 559 -44 567 44
rect 584 -44 592 44
rect 559 -50 592 -44
rect 607 44 640 50
rect 607 -44 615 44
rect 632 -44 640 44
rect 607 -50 640 -44
rect 655 44 688 50
rect 655 -44 663 44
rect 680 -44 688 44
rect 655 -50 688 -44
rect 703 44 736 50
rect 703 -44 711 44
rect 728 -44 736 44
rect 703 -50 736 -44
rect 751 44 784 50
rect 751 -44 759 44
rect 776 -44 784 44
rect 751 -50 784 -44
rect 799 44 832 50
rect 799 -44 807 44
rect 824 -44 832 44
rect 799 -50 832 -44
rect 847 44 880 50
rect 847 -44 855 44
rect 872 -44 880 44
rect 847 -50 880 -44
rect 895 44 928 50
rect 895 -44 903 44
rect 920 -44 928 44
rect 895 -50 928 -44
rect 943 44 976 50
rect 943 -44 951 44
rect 968 -44 976 44
rect 943 -50 976 -44
rect 991 44 1024 50
rect 991 -44 999 44
rect 1016 -44 1024 44
rect 991 -50 1024 -44
rect 1039 44 1072 50
rect 1039 -44 1047 44
rect 1064 -44 1072 44
rect 1039 -50 1072 -44
rect 1087 44 1120 50
rect 1087 -44 1095 44
rect 1112 -44 1120 44
rect 1087 -50 1120 -44
rect 1135 44 1168 50
rect 1135 -44 1143 44
rect 1160 -44 1168 44
rect 1135 -50 1168 -44
rect 1183 44 1216 50
rect 1183 -44 1191 44
rect 1208 -44 1216 44
rect 1183 -50 1216 -44
rect 1231 44 1264 50
rect 1231 -44 1239 44
rect 1256 -44 1264 44
rect 1231 -50 1264 -44
rect 1279 44 1312 50
rect 1279 -44 1287 44
rect 1304 -44 1312 44
rect 1279 -50 1312 -44
rect 1327 44 1360 50
rect 1327 -44 1335 44
rect 1352 -44 1360 44
rect 1327 -50 1360 -44
rect 1375 44 1408 50
rect 1375 -44 1383 44
rect 1400 -44 1408 44
rect 1375 -50 1408 -44
rect 1423 44 1454 50
rect 1423 -44 1431 44
rect 1448 -44 1454 44
rect 1423 -50 1454 -44
<< ndiffc >>
rect -1449 -44 -1432 44
rect -1401 -44 -1384 44
rect -1353 -44 -1336 44
rect -1305 -44 -1288 44
rect -1257 -44 -1240 44
rect -1209 -44 -1192 44
rect -1161 -44 -1144 44
rect -1113 -44 -1096 44
rect -1065 -44 -1048 44
rect -1017 -44 -1000 44
rect -969 -44 -952 44
rect -921 -44 -904 44
rect -873 -44 -856 44
rect -825 -44 -808 44
rect -777 -44 -760 44
rect -729 -44 -712 44
rect -681 -44 -664 44
rect -633 -44 -616 44
rect -585 -44 -568 44
rect -537 -44 -520 44
rect -489 -44 -472 44
rect -441 -44 -424 44
rect -393 -44 -376 44
rect -345 -44 -328 44
rect -297 -44 -280 44
rect -249 -44 -232 44
rect -201 -44 -184 44
rect -153 -44 -136 44
rect -105 -44 -88 44
rect -57 -44 -40 44
rect -9 -44 8 44
rect 39 -44 56 44
rect 87 -44 104 44
rect 135 -44 152 44
rect 183 -44 200 44
rect 231 -44 248 44
rect 279 -44 296 44
rect 327 -44 344 44
rect 375 -44 392 44
rect 423 -44 440 44
rect 471 -44 488 44
rect 519 -44 536 44
rect 567 -44 584 44
rect 615 -44 632 44
rect 663 -44 680 44
rect 711 -44 728 44
rect 759 -44 776 44
rect 807 -44 824 44
rect 855 -44 872 44
rect 903 -44 920 44
rect 951 -44 968 44
rect 999 -44 1016 44
rect 1047 -44 1064 44
rect 1095 -44 1112 44
rect 1143 -44 1160 44
rect 1191 -44 1208 44
rect 1239 -44 1256 44
rect 1287 -44 1304 44
rect 1335 -44 1352 44
rect 1383 -44 1400 44
rect 1431 -44 1448 44
<< psubdiff >>
rect -1506 120 -1458 137
rect 1457 120 1505 137
rect -1506 89 -1489 120
rect 1488 89 1505 120
rect -1506 -120 -1489 -89
rect 1488 -120 1505 -89
rect -1506 -137 -1458 -120
rect 1457 -137 1505 -120
<< psubdiffcont >>
rect -1458 120 1457 137
rect -1506 -89 -1489 89
rect 1488 -89 1505 89
rect -1458 -137 1457 -120
<< poly >>
rect -1424 50 -1409 63
rect -1376 50 -1361 63
rect -1328 50 -1313 63
rect -1280 50 -1265 63
rect -1232 50 -1217 63
rect -1184 50 -1169 63
rect -1136 50 -1121 63
rect -1088 50 -1073 63
rect -1040 50 -1025 63
rect -992 50 -977 63
rect -944 50 -929 63
rect -896 50 -881 63
rect -848 50 -833 63
rect -800 50 -785 63
rect -752 50 -737 63
rect -704 50 -689 63
rect -656 50 -641 63
rect -608 50 -593 63
rect -560 50 -545 63
rect -512 50 -497 63
rect -464 50 -449 63
rect -416 50 -401 63
rect -368 50 -353 63
rect -320 50 -305 63
rect -272 50 -257 63
rect -224 50 -209 63
rect -176 50 -161 63
rect -128 50 -113 63
rect -80 50 -65 63
rect -32 50 -17 63
rect 16 50 31 63
rect 64 50 79 63
rect 112 50 127 63
rect 160 50 175 63
rect 208 50 223 63
rect 256 50 271 63
rect 304 50 319 63
rect 352 50 367 63
rect 400 50 415 63
rect 448 50 463 63
rect 496 50 511 63
rect 544 50 559 63
rect 592 50 607 63
rect 640 50 655 63
rect 688 50 703 63
rect 736 50 751 63
rect 784 50 799 63
rect 832 50 847 63
rect 880 50 895 63
rect 928 50 943 63
rect 976 50 991 63
rect 1024 50 1039 63
rect 1072 50 1087 63
rect 1120 50 1135 63
rect 1168 50 1183 63
rect 1216 50 1231 63
rect 1264 50 1279 63
rect 1312 50 1327 63
rect 1360 50 1375 63
rect 1408 50 1423 63
rect -1424 -61 -1409 -50
rect -1433 -63 -1400 -61
rect -1376 -63 -1361 -50
rect -1328 -61 -1313 -50
rect -1337 -63 -1304 -61
rect -1280 -63 -1265 -50
rect -1232 -61 -1217 -50
rect -1241 -63 -1208 -61
rect -1184 -63 -1169 -50
rect -1136 -61 -1121 -50
rect -1145 -63 -1112 -61
rect -1088 -63 -1073 -50
rect -1040 -61 -1025 -50
rect -1049 -63 -1016 -61
rect -992 -63 -977 -50
rect -944 -61 -929 -50
rect -953 -63 -920 -61
rect -896 -63 -881 -50
rect -848 -61 -833 -50
rect -857 -63 -824 -61
rect -800 -63 -785 -50
rect -752 -61 -737 -50
rect -761 -63 -728 -61
rect -704 -63 -689 -50
rect -656 -61 -641 -50
rect -665 -63 -632 -61
rect -608 -63 -593 -50
rect -560 -61 -545 -50
rect -569 -63 -536 -61
rect -512 -63 -497 -50
rect -464 -61 -449 -50
rect -473 -63 -440 -61
rect -416 -63 -401 -50
rect -368 -61 -353 -50
rect -377 -63 -344 -61
rect -320 -63 -305 -50
rect -272 -61 -257 -50
rect -281 -63 -248 -61
rect -224 -63 -209 -50
rect -176 -61 -161 -50
rect -185 -63 -152 -61
rect -128 -63 -113 -50
rect -80 -61 -65 -50
rect -89 -63 -56 -61
rect -32 -63 -17 -50
rect 16 -61 31 -50
rect 7 -63 40 -61
rect 64 -63 79 -50
rect 112 -61 127 -50
rect 103 -63 136 -61
rect 160 -63 175 -50
rect 208 -61 223 -50
rect 199 -63 232 -61
rect 256 -63 271 -50
rect 304 -61 319 -50
rect 295 -63 328 -61
rect 352 -63 367 -50
rect 400 -61 415 -50
rect 391 -63 424 -61
rect 448 -63 463 -50
rect 496 -61 511 -50
rect 487 -63 520 -61
rect 544 -63 559 -50
rect 592 -61 607 -50
rect 583 -63 616 -61
rect 640 -63 655 -50
rect 688 -61 703 -50
rect 679 -63 712 -61
rect 736 -63 751 -50
rect 784 -61 799 -50
rect 775 -63 808 -61
rect 832 -63 847 -50
rect 880 -61 895 -50
rect 871 -63 904 -61
rect 928 -63 943 -50
rect 976 -61 991 -50
rect 967 -63 1000 -61
rect 1024 -63 1039 -50
rect 1072 -61 1087 -50
rect 1063 -63 1096 -61
rect 1120 -63 1135 -50
rect 1168 -61 1183 -50
rect 1159 -63 1192 -61
rect 1216 -63 1231 -50
rect 1264 -61 1279 -50
rect 1255 -63 1288 -61
rect 1312 -63 1327 -50
rect 1360 -61 1375 -50
rect 1351 -63 1384 -61
rect 1408 -63 1423 -50
rect -1433 -69 1423 -63
rect -1433 -81 -177 -69
rect -1433 -94 -1400 -81
rect -1337 -94 -1304 -81
rect -1241 -94 -1208 -81
rect -1145 -94 -1112 -81
rect -1049 -94 -1016 -81
rect -953 -94 -920 -81
rect -857 -94 -824 -81
rect -761 -94 -728 -81
rect -665 -94 -632 -81
rect -569 -94 -536 -81
rect -473 -94 -440 -81
rect -377 -94 -344 -81
rect -281 -94 -248 -81
rect -185 -86 -177 -81
rect -160 -81 1423 -69
rect -160 -86 -152 -81
rect -185 -94 -152 -86
rect -89 -94 -56 -81
rect 7 -94 40 -81
rect 103 -94 136 -81
rect 199 -94 232 -81
rect 295 -94 328 -81
rect 391 -94 424 -81
rect 487 -94 520 -81
rect 583 -94 616 -81
rect 679 -94 712 -81
rect 775 -94 808 -81
rect 871 -94 904 -81
rect 967 -94 1000 -81
rect 1063 -94 1096 -81
rect 1159 -94 1192 -81
rect 1255 -94 1288 -81
rect 1351 -94 1384 -81
<< polycont >>
rect -177 -86 -160 -69
<< locali >>
rect -1506 120 -1458 137
rect 1457 120 1505 137
rect -1506 89 -1489 120
rect 1488 89 1505 120
rect -1449 44 -1432 52
rect -1449 -52 -1432 -44
rect -1401 44 -1384 52
rect -1401 -52 -1384 -44
rect -1353 44 -1336 52
rect -1353 -52 -1336 -44
rect -1305 44 -1288 52
rect -1305 -52 -1288 -44
rect -1257 44 -1240 52
rect -1257 -52 -1240 -44
rect -1209 44 -1192 52
rect -1209 -52 -1192 -44
rect -1161 44 -1144 52
rect -1161 -52 -1144 -44
rect -1113 44 -1096 52
rect -1113 -52 -1096 -44
rect -1065 44 -1048 52
rect -1065 -52 -1048 -44
rect -1017 44 -1000 52
rect -1017 -52 -1000 -44
rect -969 44 -952 52
rect -969 -52 -952 -44
rect -921 44 -904 52
rect -921 -52 -904 -44
rect -873 44 -856 52
rect -873 -52 -856 -44
rect -825 44 -808 52
rect -825 -52 -808 -44
rect -777 44 -760 52
rect -777 -52 -760 -44
rect -729 44 -712 52
rect -729 -52 -712 -44
rect -681 44 -664 52
rect -681 -52 -664 -44
rect -633 44 -616 52
rect -633 -52 -616 -44
rect -585 44 -568 52
rect -585 -52 -568 -44
rect -537 44 -520 52
rect -537 -52 -520 -44
rect -489 44 -472 52
rect -489 -52 -472 -44
rect -441 44 -424 52
rect -441 -52 -424 -44
rect -393 44 -376 52
rect -393 -52 -376 -44
rect -345 44 -328 52
rect -345 -52 -328 -44
rect -297 44 -280 52
rect -297 -52 -280 -44
rect -249 44 -232 52
rect -249 -52 -232 -44
rect -201 44 -184 52
rect -201 -52 -184 -44
rect -153 44 -136 52
rect -153 -52 -136 -44
rect -105 44 -88 52
rect -105 -52 -88 -44
rect -57 44 -40 52
rect -57 -52 -40 -44
rect -9 44 8 52
rect -9 -52 8 -44
rect 39 44 56 52
rect 39 -52 56 -44
rect 87 44 104 52
rect 87 -52 104 -44
rect 135 44 152 52
rect 135 -52 152 -44
rect 183 44 200 52
rect 183 -52 200 -44
rect 231 44 248 52
rect 231 -52 248 -44
rect 279 44 296 52
rect 279 -52 296 -44
rect 327 44 344 52
rect 327 -52 344 -44
rect 375 44 392 52
rect 375 -52 392 -44
rect 423 44 440 52
rect 423 -52 440 -44
rect 471 44 488 52
rect 471 -52 488 -44
rect 519 44 536 52
rect 519 -52 536 -44
rect 567 44 584 52
rect 567 -52 584 -44
rect 615 44 632 52
rect 615 -52 632 -44
rect 663 44 680 52
rect 663 -52 680 -44
rect 711 44 728 52
rect 711 -52 728 -44
rect 759 44 776 52
rect 759 -52 776 -44
rect 807 44 824 52
rect 807 -52 824 -44
rect 855 44 872 52
rect 855 -52 872 -44
rect 903 44 920 52
rect 903 -52 920 -44
rect 951 44 968 52
rect 951 -52 968 -44
rect 999 44 1016 52
rect 999 -52 1016 -44
rect 1047 44 1064 52
rect 1047 -52 1064 -44
rect 1095 44 1112 52
rect 1095 -52 1112 -44
rect 1143 44 1160 52
rect 1143 -52 1160 -44
rect 1191 44 1208 52
rect 1191 -52 1208 -44
rect 1239 44 1256 52
rect 1239 -52 1256 -44
rect 1287 44 1304 52
rect 1287 -52 1304 -44
rect 1335 44 1352 52
rect 1335 -52 1352 -44
rect 1383 44 1400 52
rect 1383 -52 1400 -44
rect 1431 44 1448 52
rect 1431 -52 1448 -44
rect -185 -86 -177 -69
rect -160 -86 -152 -69
rect -1506 -120 -1489 -89
rect 1488 -120 1505 -89
rect -1506 -137 -1458 -120
rect 1457 -137 1505 -120
<< viali >>
rect -1449 -44 -1432 44
rect -1401 -44 -1384 44
rect -1353 -44 -1336 44
rect -1305 -44 -1288 44
rect -1257 -44 -1240 44
rect -1209 -44 -1192 44
rect -1161 -44 -1144 44
rect -1113 -44 -1096 44
rect -1065 -44 -1048 44
rect -1017 -44 -1000 44
rect -969 -44 -952 44
rect -921 -44 -904 44
rect -873 -44 -856 44
rect -825 -44 -808 44
rect -777 -44 -760 44
rect -729 -44 -712 44
rect -681 -44 -664 44
rect -633 -44 -616 44
rect -585 -44 -568 44
rect -537 -44 -520 44
rect -489 -44 -472 44
rect -441 -44 -424 44
rect -393 -44 -376 44
rect -345 -44 -328 44
rect -297 -44 -280 44
rect -249 -44 -232 44
rect -201 -44 -184 44
rect -153 -44 -136 44
rect -105 -44 -88 44
rect -57 -44 -40 44
rect -9 -44 8 44
rect 39 -44 56 44
rect 87 -44 104 44
rect 135 -44 152 44
rect 183 -44 200 44
rect 231 -44 248 44
rect 279 -44 296 44
rect 327 -44 344 44
rect 375 -44 392 44
rect 423 -44 440 44
rect 471 -44 488 44
rect 519 -44 536 44
rect 567 -44 584 44
rect 615 -44 632 44
rect 663 -44 680 44
rect 711 -44 728 44
rect 759 -44 776 44
rect 807 -44 824 44
rect 855 -44 872 44
rect 903 -44 920 44
rect 951 -44 968 44
rect 999 -44 1016 44
rect 1047 -44 1064 44
rect 1095 -44 1112 44
rect 1143 -44 1160 44
rect 1191 -44 1208 44
rect 1239 -44 1256 44
rect 1287 -44 1304 44
rect 1335 -44 1352 44
rect 1383 -44 1400 44
rect 1431 -44 1448 44
rect -177 -86 -160 -69
<< metal1 >>
rect -1452 44 -1429 50
rect -1452 -17 -1449 44
rect -1457 -20 -1449 -17
rect -1432 -17 -1429 44
rect -1409 47 -1376 50
rect -1409 20 -1406 47
rect -1379 20 -1376 47
rect -1409 17 -1401 20
rect -1432 -20 -1424 -17
rect -1457 -47 -1454 -20
rect -1427 -47 -1424 -20
rect -1457 -50 -1424 -47
rect -1404 -44 -1401 17
rect -1384 17 -1376 20
rect -1356 44 -1333 50
rect -1384 -44 -1381 17
rect -1356 -17 -1353 44
rect -1404 -50 -1381 -44
rect -1361 -20 -1353 -17
rect -1336 -17 -1333 44
rect -1313 47 -1280 50
rect -1313 20 -1310 47
rect -1283 20 -1280 47
rect -1313 17 -1305 20
rect -1336 -20 -1328 -17
rect -1361 -47 -1358 -20
rect -1331 -47 -1328 -20
rect -1361 -50 -1328 -47
rect -1308 -44 -1305 17
rect -1288 17 -1280 20
rect -1260 44 -1237 50
rect -1288 -44 -1285 17
rect -1260 -17 -1257 44
rect -1308 -50 -1285 -44
rect -1265 -20 -1257 -17
rect -1240 -17 -1237 44
rect -1217 47 -1184 50
rect -1217 20 -1214 47
rect -1187 20 -1184 47
rect -1217 17 -1209 20
rect -1240 -20 -1232 -17
rect -1265 -47 -1262 -20
rect -1235 -47 -1232 -20
rect -1265 -50 -1232 -47
rect -1212 -44 -1209 17
rect -1192 17 -1184 20
rect -1164 44 -1141 50
rect -1192 -44 -1189 17
rect -1164 -17 -1161 44
rect -1212 -50 -1189 -44
rect -1169 -20 -1161 -17
rect -1144 -17 -1141 44
rect -1121 47 -1088 50
rect -1121 20 -1118 47
rect -1091 20 -1088 47
rect -1121 17 -1113 20
rect -1144 -20 -1136 -17
rect -1169 -47 -1166 -20
rect -1139 -47 -1136 -20
rect -1169 -50 -1136 -47
rect -1116 -44 -1113 17
rect -1096 17 -1088 20
rect -1068 44 -1045 50
rect -1096 -44 -1093 17
rect -1068 -17 -1065 44
rect -1116 -50 -1093 -44
rect -1073 -20 -1065 -17
rect -1048 -17 -1045 44
rect -1025 47 -992 50
rect -1025 20 -1022 47
rect -995 20 -992 47
rect -1025 17 -1017 20
rect -1048 -20 -1040 -17
rect -1073 -47 -1070 -20
rect -1043 -47 -1040 -20
rect -1073 -50 -1040 -47
rect -1020 -44 -1017 17
rect -1000 17 -992 20
rect -972 44 -949 50
rect -1000 -44 -997 17
rect -972 -17 -969 44
rect -1020 -50 -997 -44
rect -977 -20 -969 -17
rect -952 -17 -949 44
rect -929 47 -896 50
rect -929 20 -926 47
rect -899 20 -896 47
rect -929 17 -921 20
rect -952 -20 -944 -17
rect -977 -47 -974 -20
rect -947 -47 -944 -20
rect -977 -50 -944 -47
rect -924 -44 -921 17
rect -904 17 -896 20
rect -876 44 -853 50
rect -904 -44 -901 17
rect -876 -17 -873 44
rect -924 -50 -901 -44
rect -881 -20 -873 -17
rect -856 -17 -853 44
rect -833 47 -800 50
rect -833 20 -830 47
rect -803 20 -800 47
rect -833 17 -825 20
rect -856 -20 -848 -17
rect -881 -47 -878 -20
rect -851 -47 -848 -20
rect -881 -50 -848 -47
rect -828 -44 -825 17
rect -808 17 -800 20
rect -780 44 -757 50
rect -808 -44 -805 17
rect -780 -17 -777 44
rect -828 -50 -805 -44
rect -785 -20 -777 -17
rect -760 -17 -757 44
rect -737 47 -704 50
rect -737 20 -734 47
rect -707 20 -704 47
rect -737 17 -729 20
rect -760 -20 -752 -17
rect -785 -47 -782 -20
rect -755 -47 -752 -20
rect -785 -50 -752 -47
rect -732 -44 -729 17
rect -712 17 -704 20
rect -684 44 -661 50
rect -712 -44 -709 17
rect -684 -17 -681 44
rect -732 -50 -709 -44
rect -689 -20 -681 -17
rect -664 -17 -661 44
rect -641 47 -608 50
rect -641 20 -638 47
rect -611 20 -608 47
rect -641 17 -633 20
rect -664 -20 -656 -17
rect -689 -47 -686 -20
rect -659 -47 -656 -20
rect -689 -50 -656 -47
rect -636 -44 -633 17
rect -616 17 -608 20
rect -588 44 -565 50
rect -616 -44 -613 17
rect -588 -17 -585 44
rect -636 -50 -613 -44
rect -593 -20 -585 -17
rect -568 -17 -565 44
rect -545 47 -512 50
rect -545 20 -542 47
rect -515 20 -512 47
rect -545 17 -537 20
rect -568 -20 -560 -17
rect -593 -47 -590 -20
rect -563 -47 -560 -20
rect -593 -50 -560 -47
rect -540 -44 -537 17
rect -520 17 -512 20
rect -492 44 -469 50
rect -520 -44 -517 17
rect -492 -17 -489 44
rect -540 -50 -517 -44
rect -497 -20 -489 -17
rect -472 -17 -469 44
rect -449 47 -416 50
rect -449 20 -446 47
rect -419 20 -416 47
rect -449 17 -441 20
rect -472 -20 -464 -17
rect -497 -47 -494 -20
rect -467 -47 -464 -20
rect -497 -50 -464 -47
rect -444 -44 -441 17
rect -424 17 -416 20
rect -396 44 -373 50
rect -424 -44 -421 17
rect -396 -17 -393 44
rect -444 -50 -421 -44
rect -401 -20 -393 -17
rect -376 -17 -373 44
rect -353 47 -320 50
rect -353 20 -350 47
rect -323 20 -320 47
rect -353 17 -345 20
rect -376 -20 -368 -17
rect -401 -47 -398 -20
rect -371 -47 -368 -20
rect -401 -50 -368 -47
rect -348 -44 -345 17
rect -328 17 -320 20
rect -300 44 -277 50
rect -328 -44 -325 17
rect -300 -17 -297 44
rect -348 -50 -325 -44
rect -305 -20 -297 -17
rect -280 -17 -277 44
rect -257 47 -224 50
rect -257 20 -254 47
rect -227 20 -224 47
rect -257 17 -249 20
rect -280 -20 -272 -17
rect -305 -47 -302 -20
rect -275 -47 -272 -20
rect -305 -50 -272 -47
rect -252 -44 -249 17
rect -232 17 -224 20
rect -204 44 -181 50
rect -232 -44 -229 17
rect -204 -17 -201 44
rect -252 -50 -229 -44
rect -209 -20 -201 -17
rect -184 -17 -181 44
rect -161 47 -128 50
rect -161 20 -158 47
rect -131 20 -128 47
rect -161 17 -153 20
rect -184 -20 -176 -17
rect -209 -47 -206 -20
rect -179 -47 -176 -20
rect -209 -50 -176 -47
rect -156 -44 -153 17
rect -136 17 -128 20
rect -108 44 -85 50
rect -136 -44 -133 17
rect -108 -17 -105 44
rect -156 -50 -133 -44
rect -113 -20 -105 -17
rect -88 -17 -85 44
rect -65 47 -32 50
rect -65 20 -62 47
rect -35 20 -32 47
rect -65 17 -57 20
rect -88 -20 -80 -17
rect -113 -47 -110 -20
rect -83 -47 -80 -20
rect -113 -50 -80 -47
rect -60 -44 -57 17
rect -40 17 -32 20
rect -12 44 11 50
rect -40 -44 -37 17
rect -12 -17 -9 44
rect -60 -50 -37 -44
rect -17 -20 -9 -17
rect 8 -17 11 44
rect 31 47 64 50
rect 31 20 34 47
rect 61 20 64 47
rect 31 17 39 20
rect 8 -20 16 -17
rect -17 -47 -14 -20
rect 13 -47 16 -20
rect -17 -50 16 -47
rect 36 -44 39 17
rect 56 17 64 20
rect 84 44 107 50
rect 56 -44 59 17
rect 84 -17 87 44
rect 36 -50 59 -44
rect 79 -20 87 -17
rect 104 -17 107 44
rect 127 47 160 50
rect 127 20 130 47
rect 157 20 160 47
rect 127 17 135 20
rect 104 -20 112 -17
rect 79 -47 82 -20
rect 109 -47 112 -20
rect 79 -50 112 -47
rect 132 -44 135 17
rect 152 17 160 20
rect 180 44 203 50
rect 152 -44 155 17
rect 180 -17 183 44
rect 132 -50 155 -44
rect 175 -20 183 -17
rect 200 -17 203 44
rect 223 47 256 50
rect 223 20 226 47
rect 253 20 256 47
rect 223 17 231 20
rect 200 -20 208 -17
rect 175 -47 178 -20
rect 205 -47 208 -20
rect 175 -50 208 -47
rect 228 -44 231 17
rect 248 17 256 20
rect 276 44 299 50
rect 248 -44 251 17
rect 276 -17 279 44
rect 228 -50 251 -44
rect 271 -20 279 -17
rect 296 -17 299 44
rect 319 47 352 50
rect 319 20 322 47
rect 349 20 352 47
rect 319 17 327 20
rect 296 -20 304 -17
rect 271 -47 274 -20
rect 301 -47 304 -20
rect 271 -50 304 -47
rect 324 -44 327 17
rect 344 17 352 20
rect 372 44 395 50
rect 344 -44 347 17
rect 372 -17 375 44
rect 324 -50 347 -44
rect 367 -20 375 -17
rect 392 -17 395 44
rect 415 47 448 50
rect 415 20 418 47
rect 445 20 448 47
rect 415 17 423 20
rect 392 -20 400 -17
rect 367 -47 370 -20
rect 397 -47 400 -20
rect 367 -50 400 -47
rect 420 -44 423 17
rect 440 17 448 20
rect 468 44 491 50
rect 440 -44 443 17
rect 468 -17 471 44
rect 420 -50 443 -44
rect 463 -20 471 -17
rect 488 -17 491 44
rect 511 47 544 50
rect 511 20 514 47
rect 541 20 544 47
rect 511 17 519 20
rect 488 -20 496 -17
rect 463 -47 466 -20
rect 493 -47 496 -20
rect 463 -50 496 -47
rect 516 -44 519 17
rect 536 17 544 20
rect 564 44 587 50
rect 536 -44 539 17
rect 564 -17 567 44
rect 516 -50 539 -44
rect 559 -20 567 -17
rect 584 -17 587 44
rect 607 47 640 50
rect 607 20 610 47
rect 637 20 640 47
rect 607 17 615 20
rect 584 -20 592 -17
rect 559 -47 562 -20
rect 589 -47 592 -20
rect 559 -50 592 -47
rect 612 -44 615 17
rect 632 17 640 20
rect 660 44 683 50
rect 632 -44 635 17
rect 660 -17 663 44
rect 612 -50 635 -44
rect 655 -20 663 -17
rect 680 -17 683 44
rect 703 47 736 50
rect 703 20 706 47
rect 733 20 736 47
rect 703 17 711 20
rect 680 -20 688 -17
rect 655 -47 658 -20
rect 685 -47 688 -20
rect 655 -50 688 -47
rect 708 -44 711 17
rect 728 17 736 20
rect 756 44 779 50
rect 728 -44 731 17
rect 756 -17 759 44
rect 708 -50 731 -44
rect 751 -20 759 -17
rect 776 -17 779 44
rect 799 47 832 50
rect 799 20 802 47
rect 829 20 832 47
rect 799 17 807 20
rect 776 -20 784 -17
rect 751 -47 754 -20
rect 781 -47 784 -20
rect 751 -50 784 -47
rect 804 -44 807 17
rect 824 17 832 20
rect 852 44 875 50
rect 824 -44 827 17
rect 852 -17 855 44
rect 804 -50 827 -44
rect 847 -20 855 -17
rect 872 -17 875 44
rect 895 47 928 50
rect 895 20 898 47
rect 925 20 928 47
rect 895 17 903 20
rect 872 -20 880 -17
rect 847 -47 850 -20
rect 877 -47 880 -20
rect 847 -50 880 -47
rect 900 -44 903 17
rect 920 17 928 20
rect 948 44 971 50
rect 920 -44 923 17
rect 948 -17 951 44
rect 900 -50 923 -44
rect 943 -20 951 -17
rect 968 -17 971 44
rect 991 47 1024 50
rect 991 20 994 47
rect 1021 20 1024 47
rect 991 17 999 20
rect 968 -20 976 -17
rect 943 -47 946 -20
rect 973 -47 976 -20
rect 943 -50 976 -47
rect 996 -44 999 17
rect 1016 17 1024 20
rect 1044 44 1067 50
rect 1016 -44 1019 17
rect 1044 -17 1047 44
rect 996 -50 1019 -44
rect 1039 -20 1047 -17
rect 1064 -17 1067 44
rect 1087 47 1120 50
rect 1087 20 1090 47
rect 1117 20 1120 47
rect 1087 17 1095 20
rect 1064 -20 1072 -17
rect 1039 -47 1042 -20
rect 1069 -47 1072 -20
rect 1039 -50 1072 -47
rect 1092 -44 1095 17
rect 1112 17 1120 20
rect 1140 44 1163 50
rect 1112 -44 1115 17
rect 1140 -17 1143 44
rect 1092 -50 1115 -44
rect 1135 -20 1143 -17
rect 1160 -17 1163 44
rect 1183 47 1216 50
rect 1183 20 1186 47
rect 1213 20 1216 47
rect 1183 17 1191 20
rect 1160 -20 1168 -17
rect 1135 -47 1138 -20
rect 1165 -47 1168 -20
rect 1135 -50 1168 -47
rect 1188 -44 1191 17
rect 1208 17 1216 20
rect 1236 44 1259 50
rect 1208 -44 1211 17
rect 1236 -17 1239 44
rect 1188 -50 1211 -44
rect 1231 -20 1239 -17
rect 1256 -17 1259 44
rect 1279 47 1312 50
rect 1279 20 1282 47
rect 1309 20 1312 47
rect 1279 17 1287 20
rect 1256 -20 1264 -17
rect 1231 -47 1234 -20
rect 1261 -47 1264 -20
rect 1231 -50 1264 -47
rect 1284 -44 1287 17
rect 1304 17 1312 20
rect 1332 44 1355 50
rect 1304 -44 1307 17
rect 1332 -17 1335 44
rect 1284 -50 1307 -44
rect 1327 -20 1335 -17
rect 1352 -17 1355 44
rect 1375 47 1408 50
rect 1375 20 1378 47
rect 1405 20 1408 47
rect 1375 17 1383 20
rect 1352 -20 1360 -17
rect 1327 -47 1330 -20
rect 1357 -47 1360 -20
rect 1327 -50 1360 -47
rect 1380 -44 1383 17
rect 1400 17 1408 20
rect 1428 44 1451 50
rect 1400 -44 1403 17
rect 1428 -17 1431 44
rect 1380 -50 1403 -44
rect 1423 -20 1431 -17
rect 1448 -17 1451 44
rect 1448 -20 1456 -17
rect 1423 -47 1426 -20
rect 1453 -47 1456 -20
rect 1423 -50 1456 -47
rect -1433 -69 1423 -66
rect -1433 -86 -177 -69
rect -160 -86 1423 -69
rect -1433 -89 1423 -86
<< via1 >>
rect -1406 44 -1379 47
rect -1406 20 -1401 44
rect -1401 20 -1384 44
rect -1384 20 -1379 44
rect -1454 -44 -1449 -20
rect -1449 -44 -1432 -20
rect -1432 -44 -1427 -20
rect -1454 -47 -1427 -44
rect -1310 44 -1283 47
rect -1310 20 -1305 44
rect -1305 20 -1288 44
rect -1288 20 -1283 44
rect -1358 -44 -1353 -20
rect -1353 -44 -1336 -20
rect -1336 -44 -1331 -20
rect -1358 -47 -1331 -44
rect -1214 44 -1187 47
rect -1214 20 -1209 44
rect -1209 20 -1192 44
rect -1192 20 -1187 44
rect -1262 -44 -1257 -20
rect -1257 -44 -1240 -20
rect -1240 -44 -1235 -20
rect -1262 -47 -1235 -44
rect -1118 44 -1091 47
rect -1118 20 -1113 44
rect -1113 20 -1096 44
rect -1096 20 -1091 44
rect -1166 -44 -1161 -20
rect -1161 -44 -1144 -20
rect -1144 -44 -1139 -20
rect -1166 -47 -1139 -44
rect -1022 44 -995 47
rect -1022 20 -1017 44
rect -1017 20 -1000 44
rect -1000 20 -995 44
rect -1070 -44 -1065 -20
rect -1065 -44 -1048 -20
rect -1048 -44 -1043 -20
rect -1070 -47 -1043 -44
rect -926 44 -899 47
rect -926 20 -921 44
rect -921 20 -904 44
rect -904 20 -899 44
rect -974 -44 -969 -20
rect -969 -44 -952 -20
rect -952 -44 -947 -20
rect -974 -47 -947 -44
rect -830 44 -803 47
rect -830 20 -825 44
rect -825 20 -808 44
rect -808 20 -803 44
rect -878 -44 -873 -20
rect -873 -44 -856 -20
rect -856 -44 -851 -20
rect -878 -47 -851 -44
rect -734 44 -707 47
rect -734 20 -729 44
rect -729 20 -712 44
rect -712 20 -707 44
rect -782 -44 -777 -20
rect -777 -44 -760 -20
rect -760 -44 -755 -20
rect -782 -47 -755 -44
rect -638 44 -611 47
rect -638 20 -633 44
rect -633 20 -616 44
rect -616 20 -611 44
rect -686 -44 -681 -20
rect -681 -44 -664 -20
rect -664 -44 -659 -20
rect -686 -47 -659 -44
rect -542 44 -515 47
rect -542 20 -537 44
rect -537 20 -520 44
rect -520 20 -515 44
rect -590 -44 -585 -20
rect -585 -44 -568 -20
rect -568 -44 -563 -20
rect -590 -47 -563 -44
rect -446 44 -419 47
rect -446 20 -441 44
rect -441 20 -424 44
rect -424 20 -419 44
rect -494 -44 -489 -20
rect -489 -44 -472 -20
rect -472 -44 -467 -20
rect -494 -47 -467 -44
rect -350 44 -323 47
rect -350 20 -345 44
rect -345 20 -328 44
rect -328 20 -323 44
rect -398 -44 -393 -20
rect -393 -44 -376 -20
rect -376 -44 -371 -20
rect -398 -47 -371 -44
rect -254 44 -227 47
rect -254 20 -249 44
rect -249 20 -232 44
rect -232 20 -227 44
rect -302 -44 -297 -20
rect -297 -44 -280 -20
rect -280 -44 -275 -20
rect -302 -47 -275 -44
rect -158 44 -131 47
rect -158 20 -153 44
rect -153 20 -136 44
rect -136 20 -131 44
rect -206 -44 -201 -20
rect -201 -44 -184 -20
rect -184 -44 -179 -20
rect -206 -47 -179 -44
rect -62 44 -35 47
rect -62 20 -57 44
rect -57 20 -40 44
rect -40 20 -35 44
rect -110 -44 -105 -20
rect -105 -44 -88 -20
rect -88 -44 -83 -20
rect -110 -47 -83 -44
rect 34 44 61 47
rect 34 20 39 44
rect 39 20 56 44
rect 56 20 61 44
rect -14 -44 -9 -20
rect -9 -44 8 -20
rect 8 -44 13 -20
rect -14 -47 13 -44
rect 130 44 157 47
rect 130 20 135 44
rect 135 20 152 44
rect 152 20 157 44
rect 82 -44 87 -20
rect 87 -44 104 -20
rect 104 -44 109 -20
rect 82 -47 109 -44
rect 226 44 253 47
rect 226 20 231 44
rect 231 20 248 44
rect 248 20 253 44
rect 178 -44 183 -20
rect 183 -44 200 -20
rect 200 -44 205 -20
rect 178 -47 205 -44
rect 322 44 349 47
rect 322 20 327 44
rect 327 20 344 44
rect 344 20 349 44
rect 274 -44 279 -20
rect 279 -44 296 -20
rect 296 -44 301 -20
rect 274 -47 301 -44
rect 418 44 445 47
rect 418 20 423 44
rect 423 20 440 44
rect 440 20 445 44
rect 370 -44 375 -20
rect 375 -44 392 -20
rect 392 -44 397 -20
rect 370 -47 397 -44
rect 514 44 541 47
rect 514 20 519 44
rect 519 20 536 44
rect 536 20 541 44
rect 466 -44 471 -20
rect 471 -44 488 -20
rect 488 -44 493 -20
rect 466 -47 493 -44
rect 610 44 637 47
rect 610 20 615 44
rect 615 20 632 44
rect 632 20 637 44
rect 562 -44 567 -20
rect 567 -44 584 -20
rect 584 -44 589 -20
rect 562 -47 589 -44
rect 706 44 733 47
rect 706 20 711 44
rect 711 20 728 44
rect 728 20 733 44
rect 658 -44 663 -20
rect 663 -44 680 -20
rect 680 -44 685 -20
rect 658 -47 685 -44
rect 802 44 829 47
rect 802 20 807 44
rect 807 20 824 44
rect 824 20 829 44
rect 754 -44 759 -20
rect 759 -44 776 -20
rect 776 -44 781 -20
rect 754 -47 781 -44
rect 898 44 925 47
rect 898 20 903 44
rect 903 20 920 44
rect 920 20 925 44
rect 850 -44 855 -20
rect 855 -44 872 -20
rect 872 -44 877 -20
rect 850 -47 877 -44
rect 994 44 1021 47
rect 994 20 999 44
rect 999 20 1016 44
rect 1016 20 1021 44
rect 946 -44 951 -20
rect 951 -44 968 -20
rect 968 -44 973 -20
rect 946 -47 973 -44
rect 1090 44 1117 47
rect 1090 20 1095 44
rect 1095 20 1112 44
rect 1112 20 1117 44
rect 1042 -44 1047 -20
rect 1047 -44 1064 -20
rect 1064 -44 1069 -20
rect 1042 -47 1069 -44
rect 1186 44 1213 47
rect 1186 20 1191 44
rect 1191 20 1208 44
rect 1208 20 1213 44
rect 1138 -44 1143 -20
rect 1143 -44 1160 -20
rect 1160 -44 1165 -20
rect 1138 -47 1165 -44
rect 1282 44 1309 47
rect 1282 20 1287 44
rect 1287 20 1304 44
rect 1304 20 1309 44
rect 1234 -44 1239 -20
rect 1239 -44 1256 -20
rect 1256 -44 1261 -20
rect 1234 -47 1261 -44
rect 1378 44 1405 47
rect 1378 20 1383 44
rect 1383 20 1400 44
rect 1400 20 1405 44
rect 1330 -44 1335 -20
rect 1335 -44 1352 -20
rect 1352 -44 1357 -20
rect 1330 -47 1357 -44
rect 1426 -44 1431 -20
rect 1431 -44 1448 -20
rect 1448 -44 1453 -20
rect 1426 -47 1453 -44
<< metal2 >>
rect -1457 47 1458 94
rect -1457 20 -1406 47
rect -1379 20 -1310 47
rect -1283 20 -1214 47
rect -1187 20 -1118 47
rect -1091 20 -1022 47
rect -995 20 -926 47
rect -899 20 -830 47
rect -803 20 -734 47
rect -707 20 -638 47
rect -611 20 -542 47
rect -515 20 -446 47
rect -419 20 -350 47
rect -323 20 -254 47
rect -227 20 -158 47
rect -131 20 -62 47
rect -35 20 34 47
rect 61 20 130 47
rect 157 20 226 47
rect 253 20 322 47
rect 349 20 418 47
rect 445 20 514 47
rect 541 20 610 47
rect 637 20 706 47
rect 733 20 802 47
rect 829 20 898 47
rect 925 20 994 47
rect 1021 20 1090 47
rect 1117 20 1186 47
rect 1213 20 1282 47
rect 1309 20 1378 47
rect 1405 20 1458 47
rect -1457 17 1458 20
rect -1457 -20 1458 -17
rect -1457 -47 -1454 -20
rect -1427 -47 -1358 -20
rect -1331 -47 -1262 -20
rect -1235 -47 -1166 -20
rect -1139 -47 -1070 -20
rect -1043 -47 -974 -20
rect -947 -47 -878 -20
rect -851 -47 -782 -20
rect -755 -47 -686 -20
rect -659 -47 -590 -20
rect -563 -47 -494 -20
rect -467 -47 -398 -20
rect -371 -47 -302 -20
rect -275 -47 -206 -20
rect -179 -47 -110 -20
rect -83 -47 -14 -20
rect 13 -47 82 -20
rect 109 -47 178 -20
rect 205 -47 274 -20
rect 301 -47 370 -20
rect 397 -47 466 -20
rect 493 -47 562 -20
rect 589 -47 658 -20
rect 685 -47 754 -20
rect 781 -47 850 -20
rect 877 -47 946 -20
rect 973 -47 1042 -20
rect 1069 -47 1138 -20
rect 1165 -47 1234 -20
rect 1261 -47 1330 -20
rect 1357 -47 1426 -20
rect 1453 -47 1458 -20
rect -1457 -94 1458 -47
<< properties >>
string FIXED_BBOX -1497 -128 1497 128
string gencell sky130_fd_pr__nfet_01v8_lvt
string library sky130
string parameters w 1.0 l 0.15 m 1 nf 60 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
