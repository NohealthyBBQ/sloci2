magic
tech sky130A
magscale 1 2
timestamp 1671759029
<< nwell >>
rect -3831 -1019 3831 1019
<< pmoslvt >>
rect -3635 -800 -3235 800
rect -3177 -800 -2777 800
rect -2719 -800 -2319 800
rect -2261 -800 -1861 800
rect -1803 -800 -1403 800
rect -1345 -800 -945 800
rect -887 -800 -487 800
rect -429 -800 -29 800
rect 29 -800 429 800
rect 487 -800 887 800
rect 945 -800 1345 800
rect 1403 -800 1803 800
rect 1861 -800 2261 800
rect 2319 -800 2719 800
rect 2777 -800 3177 800
rect 3235 -800 3635 800
<< pdiff >>
rect -3693 788 -3635 800
rect -3693 -788 -3681 788
rect -3647 -788 -3635 788
rect -3693 -800 -3635 -788
rect -3235 788 -3177 800
rect -3235 -788 -3223 788
rect -3189 -788 -3177 788
rect -3235 -800 -3177 -788
rect -2777 788 -2719 800
rect -2777 -788 -2765 788
rect -2731 -788 -2719 788
rect -2777 -800 -2719 -788
rect -2319 788 -2261 800
rect -2319 -788 -2307 788
rect -2273 -788 -2261 788
rect -2319 -800 -2261 -788
rect -1861 788 -1803 800
rect -1861 -788 -1849 788
rect -1815 -788 -1803 788
rect -1861 -800 -1803 -788
rect -1403 788 -1345 800
rect -1403 -788 -1391 788
rect -1357 -788 -1345 788
rect -1403 -800 -1345 -788
rect -945 788 -887 800
rect -945 -788 -933 788
rect -899 -788 -887 788
rect -945 -800 -887 -788
rect -487 788 -429 800
rect -487 -788 -475 788
rect -441 -788 -429 788
rect -487 -800 -429 -788
rect -29 788 29 800
rect -29 -788 -17 788
rect 17 -788 29 788
rect -29 -800 29 -788
rect 429 788 487 800
rect 429 -788 441 788
rect 475 -788 487 788
rect 429 -800 487 -788
rect 887 788 945 800
rect 887 -788 899 788
rect 933 -788 945 788
rect 887 -800 945 -788
rect 1345 788 1403 800
rect 1345 -788 1357 788
rect 1391 -788 1403 788
rect 1345 -800 1403 -788
rect 1803 788 1861 800
rect 1803 -788 1815 788
rect 1849 -788 1861 788
rect 1803 -800 1861 -788
rect 2261 788 2319 800
rect 2261 -788 2273 788
rect 2307 -788 2319 788
rect 2261 -800 2319 -788
rect 2719 788 2777 800
rect 2719 -788 2731 788
rect 2765 -788 2777 788
rect 2719 -800 2777 -788
rect 3177 788 3235 800
rect 3177 -788 3189 788
rect 3223 -788 3235 788
rect 3177 -800 3235 -788
rect 3635 788 3693 800
rect 3635 -788 3647 788
rect 3681 -788 3693 788
rect 3635 -800 3693 -788
<< pdiffc >>
rect -3681 -788 -3647 788
rect -3223 -788 -3189 788
rect -2765 -788 -2731 788
rect -2307 -788 -2273 788
rect -1849 -788 -1815 788
rect -1391 -788 -1357 788
rect -933 -788 -899 788
rect -475 -788 -441 788
rect -17 -788 17 788
rect 441 -788 475 788
rect 899 -788 933 788
rect 1357 -788 1391 788
rect 1815 -788 1849 788
rect 2273 -788 2307 788
rect 2731 -788 2765 788
rect 3189 -788 3223 788
rect 3647 -788 3681 788
<< nsubdiff >>
rect -3795 949 3795 983
rect -3795 887 -3761 949
rect 3761 887 3795 949
rect -3795 -949 -3761 -887
rect 3761 -949 3795 -887
rect -3795 -983 3795 -949
<< nsubdiffcont >>
rect -3795 -887 -3761 887
rect 3761 -887 3795 887
<< poly >>
rect -3635 881 -3235 897
rect -3635 847 -3619 881
rect -3251 847 -3235 881
rect -3635 800 -3235 847
rect -3177 881 -2777 897
rect -3177 847 -3161 881
rect -2793 847 -2777 881
rect -3177 800 -2777 847
rect -2719 881 -2319 897
rect -2719 847 -2703 881
rect -2335 847 -2319 881
rect -2719 800 -2319 847
rect -2261 881 -1861 897
rect -2261 847 -2245 881
rect -1877 847 -1861 881
rect -2261 800 -1861 847
rect -1803 881 -1403 897
rect -1803 847 -1787 881
rect -1419 847 -1403 881
rect -1803 800 -1403 847
rect -1345 881 -945 897
rect -1345 847 -1329 881
rect -961 847 -945 881
rect -1345 800 -945 847
rect -887 881 -487 897
rect -887 847 -871 881
rect -503 847 -487 881
rect -887 800 -487 847
rect -429 881 -29 897
rect -429 847 -413 881
rect -45 847 -29 881
rect -429 800 -29 847
rect 29 881 429 897
rect 29 847 45 881
rect 413 847 429 881
rect 29 800 429 847
rect 487 881 887 897
rect 487 847 503 881
rect 871 847 887 881
rect 487 800 887 847
rect 945 881 1345 897
rect 945 847 961 881
rect 1329 847 1345 881
rect 945 800 1345 847
rect 1403 881 1803 897
rect 1403 847 1419 881
rect 1787 847 1803 881
rect 1403 800 1803 847
rect 1861 881 2261 897
rect 1861 847 1877 881
rect 2245 847 2261 881
rect 1861 800 2261 847
rect 2319 881 2719 897
rect 2319 847 2335 881
rect 2703 847 2719 881
rect 2319 800 2719 847
rect 2777 881 3177 897
rect 2777 847 2793 881
rect 3161 847 3177 881
rect 2777 800 3177 847
rect 3235 881 3635 897
rect 3235 847 3251 881
rect 3619 847 3635 881
rect 3235 800 3635 847
rect -3635 -847 -3235 -800
rect -3635 -881 -3619 -847
rect -3251 -881 -3235 -847
rect -3635 -897 -3235 -881
rect -3177 -847 -2777 -800
rect -3177 -881 -3161 -847
rect -2793 -881 -2777 -847
rect -3177 -897 -2777 -881
rect -2719 -847 -2319 -800
rect -2719 -881 -2703 -847
rect -2335 -881 -2319 -847
rect -2719 -897 -2319 -881
rect -2261 -847 -1861 -800
rect -2261 -881 -2245 -847
rect -1877 -881 -1861 -847
rect -2261 -897 -1861 -881
rect -1803 -847 -1403 -800
rect -1803 -881 -1787 -847
rect -1419 -881 -1403 -847
rect -1803 -897 -1403 -881
rect -1345 -847 -945 -800
rect -1345 -881 -1329 -847
rect -961 -881 -945 -847
rect -1345 -897 -945 -881
rect -887 -847 -487 -800
rect -887 -881 -871 -847
rect -503 -881 -487 -847
rect -887 -897 -487 -881
rect -429 -847 -29 -800
rect -429 -881 -413 -847
rect -45 -881 -29 -847
rect -429 -897 -29 -881
rect 29 -847 429 -800
rect 29 -881 45 -847
rect 413 -881 429 -847
rect 29 -897 429 -881
rect 487 -847 887 -800
rect 487 -881 503 -847
rect 871 -881 887 -847
rect 487 -897 887 -881
rect 945 -847 1345 -800
rect 945 -881 961 -847
rect 1329 -881 1345 -847
rect 945 -897 1345 -881
rect 1403 -847 1803 -800
rect 1403 -881 1419 -847
rect 1787 -881 1803 -847
rect 1403 -897 1803 -881
rect 1861 -847 2261 -800
rect 1861 -881 1877 -847
rect 2245 -881 2261 -847
rect 1861 -897 2261 -881
rect 2319 -847 2719 -800
rect 2319 -881 2335 -847
rect 2703 -881 2719 -847
rect 2319 -897 2719 -881
rect 2777 -847 3177 -800
rect 2777 -881 2793 -847
rect 3161 -881 3177 -847
rect 2777 -897 3177 -881
rect 3235 -847 3635 -800
rect 3235 -881 3251 -847
rect 3619 -881 3635 -847
rect 3235 -897 3635 -881
<< polycont >>
rect -3619 847 -3251 881
rect -3161 847 -2793 881
rect -2703 847 -2335 881
rect -2245 847 -1877 881
rect -1787 847 -1419 881
rect -1329 847 -961 881
rect -871 847 -503 881
rect -413 847 -45 881
rect 45 847 413 881
rect 503 847 871 881
rect 961 847 1329 881
rect 1419 847 1787 881
rect 1877 847 2245 881
rect 2335 847 2703 881
rect 2793 847 3161 881
rect 3251 847 3619 881
rect -3619 -881 -3251 -847
rect -3161 -881 -2793 -847
rect -2703 -881 -2335 -847
rect -2245 -881 -1877 -847
rect -1787 -881 -1419 -847
rect -1329 -881 -961 -847
rect -871 -881 -503 -847
rect -413 -881 -45 -847
rect 45 -881 413 -847
rect 503 -881 871 -847
rect 961 -881 1329 -847
rect 1419 -881 1787 -847
rect 1877 -881 2245 -847
rect 2335 -881 2703 -847
rect 2793 -881 3161 -847
rect 3251 -881 3619 -847
<< locali >>
rect -3795 949 3795 983
rect -3795 887 -3761 949
rect 3761 887 3795 949
rect -3635 847 -3619 881
rect -3251 847 -3235 881
rect -3177 847 -3161 881
rect -2793 847 -2777 881
rect -2719 847 -2703 881
rect -2335 847 -2319 881
rect -2261 847 -2245 881
rect -1877 847 -1861 881
rect -1803 847 -1787 881
rect -1419 847 -1403 881
rect -1345 847 -1329 881
rect -961 847 -945 881
rect -887 847 -871 881
rect -503 847 -487 881
rect -429 847 -413 881
rect -45 847 -29 881
rect 29 847 45 881
rect 413 847 429 881
rect 487 847 503 881
rect 871 847 887 881
rect 945 847 961 881
rect 1329 847 1345 881
rect 1403 847 1419 881
rect 1787 847 1803 881
rect 1861 847 1877 881
rect 2245 847 2261 881
rect 2319 847 2335 881
rect 2703 847 2719 881
rect 2777 847 2793 881
rect 3161 847 3177 881
rect 3235 847 3251 881
rect 3619 847 3635 881
rect -3681 788 -3647 804
rect -3681 -804 -3647 -788
rect -3223 788 -3189 804
rect -3223 -804 -3189 -788
rect -2765 788 -2731 804
rect -2765 -804 -2731 -788
rect -2307 788 -2273 804
rect -2307 -804 -2273 -788
rect -1849 788 -1815 804
rect -1849 -804 -1815 -788
rect -1391 788 -1357 804
rect -1391 -804 -1357 -788
rect -933 788 -899 804
rect -933 -804 -899 -788
rect -475 788 -441 804
rect -475 -804 -441 -788
rect -17 788 17 804
rect -17 -804 17 -788
rect 441 788 475 804
rect 441 -804 475 -788
rect 899 788 933 804
rect 899 -804 933 -788
rect 1357 788 1391 804
rect 1357 -804 1391 -788
rect 1815 788 1849 804
rect 1815 -804 1849 -788
rect 2273 788 2307 804
rect 2273 -804 2307 -788
rect 2731 788 2765 804
rect 2731 -804 2765 -788
rect 3189 788 3223 804
rect 3189 -804 3223 -788
rect 3647 788 3681 804
rect 3647 -804 3681 -788
rect -3635 -881 -3619 -847
rect -3251 -881 -3235 -847
rect -3177 -881 -3161 -847
rect -2793 -881 -2777 -847
rect -2719 -881 -2703 -847
rect -2335 -881 -2319 -847
rect -2261 -881 -2245 -847
rect -1877 -881 -1861 -847
rect -1803 -881 -1787 -847
rect -1419 -881 -1403 -847
rect -1345 -881 -1329 -847
rect -961 -881 -945 -847
rect -887 -881 -871 -847
rect -503 -881 -487 -847
rect -429 -881 -413 -847
rect -45 -881 -29 -847
rect 29 -881 45 -847
rect 413 -881 429 -847
rect 487 -881 503 -847
rect 871 -881 887 -847
rect 945 -881 961 -847
rect 1329 -881 1345 -847
rect 1403 -881 1419 -847
rect 1787 -881 1803 -847
rect 1861 -881 1877 -847
rect 2245 -881 2261 -847
rect 2319 -881 2335 -847
rect 2703 -881 2719 -847
rect 2777 -881 2793 -847
rect 3161 -881 3177 -847
rect 3235 -881 3251 -847
rect 3619 -881 3635 -847
rect -3795 -949 -3761 -887
rect 3761 -949 3795 -887
rect -3795 -983 3795 -949
<< viali >>
rect -3619 847 -3251 881
rect -3161 847 -2793 881
rect -2703 847 -2335 881
rect -2245 847 -1877 881
rect -1787 847 -1419 881
rect -1329 847 -961 881
rect -871 847 -503 881
rect -413 847 -45 881
rect 45 847 413 881
rect 503 847 871 881
rect 961 847 1329 881
rect 1419 847 1787 881
rect 1877 847 2245 881
rect 2335 847 2703 881
rect 2793 847 3161 881
rect 3251 847 3619 881
rect -3681 -788 -3647 788
rect -3223 -788 -3189 788
rect -2765 -788 -2731 788
rect -2307 -788 -2273 788
rect -1849 -788 -1815 788
rect -1391 -788 -1357 788
rect -933 -788 -899 788
rect -475 -788 -441 788
rect -17 -788 17 788
rect 441 -788 475 788
rect 899 -788 933 788
rect 1357 -788 1391 788
rect 1815 -788 1849 788
rect 2273 -788 2307 788
rect 2731 -788 2765 788
rect 3189 -788 3223 788
rect 3647 -788 3681 788
rect -3619 -881 -3251 -847
rect -3161 -881 -2793 -847
rect -2703 -881 -2335 -847
rect -2245 -881 -1877 -847
rect -1787 -881 -1419 -847
rect -1329 -881 -961 -847
rect -871 -881 -503 -847
rect -413 -881 -45 -847
rect 45 -881 413 -847
rect 503 -881 871 -847
rect 961 -881 1329 -847
rect 1419 -881 1787 -847
rect 1877 -881 2245 -847
rect 2335 -881 2703 -847
rect 2793 -881 3161 -847
rect 3251 -881 3619 -847
<< metal1 >>
rect -3631 881 -3239 887
rect -3631 847 -3619 881
rect -3251 847 -3239 881
rect -3631 841 -3239 847
rect -3173 881 -2781 887
rect -3173 847 -3161 881
rect -2793 847 -2781 881
rect -3173 841 -2781 847
rect -2715 881 -2323 887
rect -2715 847 -2703 881
rect -2335 847 -2323 881
rect -2715 841 -2323 847
rect -2257 881 -1865 887
rect -2257 847 -2245 881
rect -1877 847 -1865 881
rect -2257 841 -1865 847
rect -1799 881 -1407 887
rect -1799 847 -1787 881
rect -1419 847 -1407 881
rect -1799 841 -1407 847
rect -1341 881 -949 887
rect -1341 847 -1329 881
rect -961 847 -949 881
rect -1341 841 -949 847
rect -883 881 -491 887
rect -883 847 -871 881
rect -503 847 -491 881
rect -883 841 -491 847
rect -425 881 -33 887
rect -425 847 -413 881
rect -45 847 -33 881
rect -425 841 -33 847
rect 33 881 425 887
rect 33 847 45 881
rect 413 847 425 881
rect 33 841 425 847
rect 491 881 883 887
rect 491 847 503 881
rect 871 847 883 881
rect 491 841 883 847
rect 949 881 1341 887
rect 949 847 961 881
rect 1329 847 1341 881
rect 949 841 1341 847
rect 1407 881 1799 887
rect 1407 847 1419 881
rect 1787 847 1799 881
rect 1407 841 1799 847
rect 1865 881 2257 887
rect 1865 847 1877 881
rect 2245 847 2257 881
rect 1865 841 2257 847
rect 2323 881 2715 887
rect 2323 847 2335 881
rect 2703 847 2715 881
rect 2323 841 2715 847
rect 2781 881 3173 887
rect 2781 847 2793 881
rect 3161 847 3173 881
rect 2781 841 3173 847
rect 3239 881 3631 887
rect 3239 847 3251 881
rect 3619 847 3631 881
rect 3239 841 3631 847
rect -3687 788 -3641 800
rect -3687 -788 -3681 788
rect -3647 -788 -3641 788
rect -3687 -800 -3641 -788
rect -3229 788 -3183 800
rect -3229 -788 -3223 788
rect -3189 -788 -3183 788
rect -3229 -800 -3183 -788
rect -2771 788 -2725 800
rect -2771 -788 -2765 788
rect -2731 -788 -2725 788
rect -2771 -800 -2725 -788
rect -2313 788 -2267 800
rect -2313 -788 -2307 788
rect -2273 -788 -2267 788
rect -2313 -800 -2267 -788
rect -1855 788 -1809 800
rect -1855 -788 -1849 788
rect -1815 -788 -1809 788
rect -1855 -800 -1809 -788
rect -1397 788 -1351 800
rect -1397 -788 -1391 788
rect -1357 -788 -1351 788
rect -1397 -800 -1351 -788
rect -939 788 -893 800
rect -939 -788 -933 788
rect -899 -788 -893 788
rect -939 -800 -893 -788
rect -481 788 -435 800
rect -481 -788 -475 788
rect -441 -788 -435 788
rect -481 -800 -435 -788
rect -23 788 23 800
rect -23 -788 -17 788
rect 17 -788 23 788
rect -23 -800 23 -788
rect 435 788 481 800
rect 435 -788 441 788
rect 475 -788 481 788
rect 435 -800 481 -788
rect 893 788 939 800
rect 893 -788 899 788
rect 933 -788 939 788
rect 893 -800 939 -788
rect 1351 788 1397 800
rect 1351 -788 1357 788
rect 1391 -788 1397 788
rect 1351 -800 1397 -788
rect 1809 788 1855 800
rect 1809 -788 1815 788
rect 1849 -788 1855 788
rect 1809 -800 1855 -788
rect 2267 788 2313 800
rect 2267 -788 2273 788
rect 2307 -788 2313 788
rect 2267 -800 2313 -788
rect 2725 788 2771 800
rect 2725 -788 2731 788
rect 2765 -788 2771 788
rect 2725 -800 2771 -788
rect 3183 788 3229 800
rect 3183 -788 3189 788
rect 3223 -788 3229 788
rect 3183 -800 3229 -788
rect 3641 788 3687 800
rect 3641 -788 3647 788
rect 3681 -788 3687 788
rect 3641 -800 3687 -788
rect -3631 -847 -3239 -841
rect -3631 -881 -3619 -847
rect -3251 -881 -3239 -847
rect -3631 -887 -3239 -881
rect -3173 -847 -2781 -841
rect -3173 -881 -3161 -847
rect -2793 -881 -2781 -847
rect -3173 -887 -2781 -881
rect -2715 -847 -2323 -841
rect -2715 -881 -2703 -847
rect -2335 -881 -2323 -847
rect -2715 -887 -2323 -881
rect -2257 -847 -1865 -841
rect -2257 -881 -2245 -847
rect -1877 -881 -1865 -847
rect -2257 -887 -1865 -881
rect -1799 -847 -1407 -841
rect -1799 -881 -1787 -847
rect -1419 -881 -1407 -847
rect -1799 -887 -1407 -881
rect -1341 -847 -949 -841
rect -1341 -881 -1329 -847
rect -961 -881 -949 -847
rect -1341 -887 -949 -881
rect -883 -847 -491 -841
rect -883 -881 -871 -847
rect -503 -881 -491 -847
rect -883 -887 -491 -881
rect -425 -847 -33 -841
rect -425 -881 -413 -847
rect -45 -881 -33 -847
rect -425 -887 -33 -881
rect 33 -847 425 -841
rect 33 -881 45 -847
rect 413 -881 425 -847
rect 33 -887 425 -881
rect 491 -847 883 -841
rect 491 -881 503 -847
rect 871 -881 883 -847
rect 491 -887 883 -881
rect 949 -847 1341 -841
rect 949 -881 961 -847
rect 1329 -881 1341 -847
rect 949 -887 1341 -881
rect 1407 -847 1799 -841
rect 1407 -881 1419 -847
rect 1787 -881 1799 -847
rect 1407 -887 1799 -881
rect 1865 -847 2257 -841
rect 1865 -881 1877 -847
rect 2245 -881 2257 -847
rect 1865 -887 2257 -881
rect 2323 -847 2715 -841
rect 2323 -881 2335 -847
rect 2703 -881 2715 -847
rect 2323 -887 2715 -881
rect 2781 -847 3173 -841
rect 2781 -881 2793 -847
rect 3161 -881 3173 -847
rect 2781 -887 3173 -881
rect 3239 -847 3631 -841
rect 3239 -881 3251 -847
rect 3619 -881 3631 -847
rect 3239 -887 3631 -881
<< properties >>
string FIXED_BBOX -3778 -966 3778 966
string gencell sky130_fd_pr__pfet_01v8_lvt
string library sky130
string parameters w 8 l 2 m 1 nf 16 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 0 gbc 0 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.35 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
