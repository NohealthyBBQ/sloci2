magic
tech sky130A
magscale 1 2
timestamp 1672523391
<< metal1 >>
rect 571790 692400 571800 692800
rect 572200 692400 572210 692800
rect 571980 691860 572060 692400
rect 571500 691780 572060 691860
rect 572590 691680 572600 691800
rect 571520 691540 572600 691680
rect 572590 691400 572600 691540
rect 573000 691400 573010 691800
rect 18200 682212 18500 682224
rect 18200 682156 18214 682212
rect 18484 682198 18500 682212
rect 18484 682156 49554 682198
rect 18200 682150 49554 682156
rect 17600 682116 17900 682128
rect 17600 682060 17614 682116
rect 17884 682102 17900 682116
rect 17884 682060 48316 682102
rect 17600 682054 48316 682060
rect 17000 682024 17300 682036
rect 17000 681968 17014 682024
rect 17284 682010 17300 682024
rect 17284 681968 47328 682010
rect 17000 681962 47328 681968
rect 16400 681932 16700 681944
rect 16400 681876 16414 681932
rect 16684 681918 16700 681932
rect 16684 681876 46008 681918
rect 16400 681870 46008 681876
rect 15800 681846 16100 681858
rect 15800 681790 15814 681846
rect 16084 681832 16100 681846
rect 45970 681832 46008 681870
rect 16084 681790 45346 681832
rect 47286 681828 47328 681962
rect 48278 681842 48316 682054
rect 49516 681820 49554 682150
rect 15800 681784 45346 681790
rect 254100 579500 254400 581700
rect 254090 578700 254100 579500
rect 254400 578700 254410 579500
rect 254100 578600 254400 578700
rect 317970 563360 317980 563420
rect 318040 563360 318050 563420
rect 309720 560380 309840 560560
rect 309720 560240 309740 560380
rect 309820 560240 309840 560380
rect 309720 560220 309840 560240
<< via1 >>
rect 571800 692400 572200 692800
rect 572600 691400 573000 691800
rect 18214 682156 18484 682212
rect 17614 682060 17884 682116
rect 17014 681968 17284 682024
rect 16414 681876 16684 681932
rect 15814 681790 16084 681846
rect 254100 578700 254400 579500
rect 317980 563360 318040 563420
rect 309740 560240 309820 560380
<< metal2 >>
rect 571800 692800 572200 692810
rect 571800 692390 572200 692400
rect 572600 691800 573000 691810
rect 572600 691390 573000 691400
rect 53000 685600 58800 685800
rect 53000 685476 57600 685600
rect 52994 685400 57600 685476
rect 58600 685400 58800 685600
rect 53000 685200 58800 685400
rect 18200 682212 18500 682224
rect 18200 682156 18214 682212
rect 18484 682156 18500 682212
rect 18200 682150 18500 682156
rect 17600 682116 17900 682128
rect 17600 682060 17614 682116
rect 17884 682060 17900 682116
rect 17600 682054 17900 682060
rect 17000 682024 17300 682036
rect 17000 681968 17014 682024
rect 17284 681968 17300 682024
rect 17000 681962 17300 681968
rect 16400 681932 16700 681944
rect 16400 681876 16414 681932
rect 16684 681876 16700 681932
rect 16400 681870 16700 681876
rect 15800 681846 16100 681858
rect 15800 681790 15814 681846
rect 16084 681790 16100 681846
rect 15800 681784 16100 681790
rect 333600 624800 334200 624810
rect 304400 624300 333600 624500
rect 304400 624100 304800 624300
rect 333600 623990 334200 624000
rect 307900 619100 308000 619110
rect 307900 618890 308000 618900
rect 311400 619100 311600 619110
rect 333900 619100 334100 619110
rect 311600 618900 333900 619100
rect 311400 618890 311600 618900
rect 333900 618890 334100 618900
rect 311500 616600 311700 616610
rect 331800 616600 332000 616610
rect 308300 616560 308380 616570
rect 308300 616450 308380 616460
rect 311700 616400 331800 616600
rect 332000 616400 332200 616600
rect 311500 616390 311700 616400
rect 331800 616390 332000 616400
rect 254100 579500 254400 579510
rect 254100 578690 254400 578700
rect 307600 566700 307800 566710
rect 307800 566500 309600 566700
rect 307600 566490 307800 566500
rect 317980 563420 318040 563430
rect 317980 563350 318040 563360
rect 309740 560380 309820 560390
rect 309740 560230 309820 560240
rect 483100 274050 565950 274200
rect 483100 273950 565500 274050
rect 565900 273950 565950 274050
rect 483100 273800 565950 273950
<< via2 >>
rect 571800 692400 572200 692800
rect 572600 691400 573000 691800
rect 57600 685400 58600 685600
rect 18214 682156 18484 682212
rect 17614 682060 17884 682116
rect 17014 681968 17284 682024
rect 16414 681876 16684 681932
rect 15814 681790 16084 681846
rect 333600 624000 334200 624800
rect 307900 618900 308000 619100
rect 311400 618900 311600 619100
rect 333900 618900 334100 619100
rect 308300 616460 308380 616560
rect 311500 616400 311700 616600
rect 331800 616400 332000 616600
rect 254100 578700 254400 579500
rect 307600 566500 307800 566700
rect 317980 563360 318040 563420
rect 309740 560240 309820 560380
rect 565500 273950 565900 274050
<< metal3 >>
rect 120194 702300 125194 704800
rect 165594 702300 170594 704800
rect 170894 702300 173094 704800
rect 173394 702300 175594 704800
rect 175894 702300 180894 704800
rect 217294 702300 222294 704800
rect 222594 702300 224794 704800
rect 225094 702300 227294 704800
rect 227594 702300 232594 704800
rect 318994 702300 323994 704800
rect 324294 702300 326494 704800
rect 326794 702300 328994 704800
rect 329294 702300 334294 704800
rect 413394 702300 418394 704800
rect 465394 702300 470394 704800
rect 510594 702340 515394 704800
rect 520594 702340 525394 704800
rect 566594 702300 571594 704800
rect 17880 690500 19240 696000
rect 69400 690500 70760 696000
rect 17880 690460 43920 690500
rect 17880 689180 43280 690460
rect 43860 689180 43920 690460
rect 17880 689140 43920 689180
rect 45740 690460 70760 690500
rect 45740 689180 45800 690460
rect 46380 689180 70760 690460
rect 45740 689140 70760 689180
rect 45004 688712 55292 688744
rect 45004 688398 54174 688712
rect 55256 688398 55292 688712
rect 45004 688346 55292 688398
rect 57590 685600 58610 685605
rect 57590 685400 57600 685600
rect 58600 685400 58610 685600
rect 57590 685395 58610 685400
rect -800 680242 1700 685242
rect 48024 682770 55292 682774
rect 44526 682700 55292 682770
rect 44526 682364 54202 682700
rect 55256 682364 55292 682700
rect 44526 682302 55292 682364
rect 44526 682298 50704 682302
rect 18200 682212 18500 682224
rect 18200 682156 18214 682212
rect 18484 682156 18500 682212
rect 17600 682116 17900 682130
rect 17600 682060 17614 682116
rect 17884 682060 17900 682116
rect 17000 682024 17300 682038
rect 17000 681968 17014 682024
rect 17284 681968 17300 682024
rect 16400 681932 16700 681946
rect 16400 681876 16414 681932
rect 16684 681876 16700 681932
rect 15800 681846 16100 681858
rect 15800 681790 15814 681846
rect 16084 681790 16100 681846
rect 5300 648680 9080 648700
rect 720 648642 9080 648680
rect -800 648570 9080 648642
rect -800 643880 5476 648570
rect -800 643842 1660 643880
rect 1818 641552 5476 643880
rect 8888 641552 9080 648570
rect -800 638640 1660 638642
rect 1818 638640 9080 641552
rect -800 638240 9080 638640
rect -800 633842 9040 638240
rect 1400 633840 9040 633842
rect 1582 564242 8000 564262
rect -800 563676 8000 564242
rect -800 559442 2434 563676
rect 1582 557958 2434 559442
rect 7216 557958 8000 563676
rect 1582 554242 8000 557958
rect -800 549442 8000 554242
rect 15800 508150 16100 681790
rect 2200 507950 16100 508150
rect 16400 464900 16700 681876
rect 2200 464700 16700 464900
rect 17000 421700 17300 681968
rect 2200 421500 17300 421700
rect 17600 378500 17900 682060
rect 2200 378300 17900 378500
rect 18200 335250 18500 682156
rect 122400 581400 123200 702300
rect 229000 654000 231000 702300
rect 569200 692800 569600 702300
rect 571790 692800 572210 692805
rect 569200 692400 571800 692800
rect 572200 692400 572210 692800
rect 571790 692395 572210 692400
rect 572590 691800 573010 691805
rect 572590 691400 572600 691800
rect 573000 691400 573010 691800
rect 572590 691395 573010 691400
rect 572600 681200 573000 691395
rect 582300 681200 584800 682984
rect 572600 680800 584800 681200
rect 582300 677984 584800 680800
rect 229000 652000 322000 654000
rect 307890 619100 308010 619105
rect 311390 619100 311610 619105
rect 307890 618900 307900 619100
rect 308000 618900 311400 619100
rect 311600 618900 311610 619100
rect 307890 618895 308010 618900
rect 311390 618895 311610 618900
rect 311490 616600 311710 616605
rect 308290 616560 308390 616565
rect 311490 616560 311500 616600
rect 308290 616460 308300 616560
rect 308380 616460 311500 616560
rect 308290 616455 308390 616460
rect 311490 616400 311500 616460
rect 311700 616400 311710 616600
rect 311490 616395 311710 616400
rect 262990 615000 263000 615800
rect 263600 615000 263610 615800
rect 260790 613400 260800 614200
rect 261400 613400 261410 614200
rect 260800 610700 261400 613400
rect 263000 610600 263600 615000
rect 293080 601240 302380 601260
rect 293080 601140 302240 601240
rect 302360 601140 302380 601240
rect 293080 601120 302380 601140
rect 293020 597720 302000 597740
rect 293020 597620 301820 597720
rect 301980 597620 302000 597720
rect 293020 597600 302000 597620
rect 122400 581200 239200 581400
rect 242700 581200 242840 583080
rect 122400 581100 242840 581200
rect 122400 581000 239200 581100
rect 254090 579500 254410 579505
rect 254090 578700 254100 579500
rect 254400 579400 254410 579500
rect 254400 578800 303400 579400
rect 254400 578700 254410 578800
rect 254090 578695 254410 578700
rect 302800 560400 303400 578800
rect 321000 567400 322000 652000
rect 582340 639784 584800 644584
rect 582340 629784 584800 634584
rect 333590 624800 334210 624805
rect 333590 624000 333600 624800
rect 334200 624000 334210 624800
rect 532790 624000 532800 624800
rect 533600 624000 533610 624800
rect 333590 623995 334210 624000
rect 333890 619100 334110 619105
rect 333890 618900 333900 619100
rect 334100 618900 334110 619100
rect 333890 618895 334110 618900
rect 331790 616600 332010 616605
rect 331790 616400 331800 616600
rect 332000 616400 332010 616600
rect 331790 616395 332010 616400
rect 307590 567000 307600 567200
rect 307800 567000 310400 567200
rect 307590 566700 307810 566705
rect 307590 566500 307600 566700
rect 307800 566500 307810 566700
rect 307590 566495 307810 566500
rect 317960 563420 318060 563440
rect 317960 563360 317980 563420
rect 318040 563360 318060 563420
rect 302800 560380 310000 560400
rect 302800 560240 309740 560380
rect 309820 560240 310000 560380
rect 302800 560200 310000 560240
rect 317960 557020 318060 563360
rect 317560 410000 318560 557020
rect 331800 453400 332000 616395
rect 333900 497800 334100 618895
rect 533000 587400 533400 624000
rect 583520 589472 584800 589584
rect 583520 588290 584800 588402
rect 533000 587220 583800 587400
rect 533000 587108 584800 587220
rect 533000 587000 583800 587108
rect 583520 585926 584800 586038
rect 583520 584744 584800 584856
rect 583520 583562 584800 583674
rect 582340 550562 584800 555362
rect 582340 540562 584800 545362
rect 583520 500050 584800 500162
rect 583520 498868 584800 498980
rect 581800 497800 583700 497900
rect 333900 497798 583700 497800
rect 333900 497686 584800 497798
rect 333900 497600 583700 497686
rect 581800 497500 583700 497600
rect 583520 496504 584800 496616
rect 583520 495322 584800 495434
rect 583520 494140 584800 494252
rect 583520 455628 584800 455740
rect 583520 454446 584800 454558
rect 582200 453400 583800 453500
rect 331800 453376 583800 453400
rect 331800 453264 584800 453376
rect 331800 453200 583800 453264
rect 582200 453100 583800 453200
rect 583520 452082 584800 452194
rect 583520 450900 584800 451012
rect 583520 449718 584800 449830
rect 583520 411206 584800 411318
rect 583520 410024 584800 410136
rect 317200 409200 581200 410000
rect 317200 408954 583800 409200
rect 317200 408842 584800 408954
rect 317200 408600 583800 408842
rect 317200 408000 581200 408600
rect 583520 407660 584800 407772
rect 583520 406478 584800 406590
rect 583520 405296 584800 405408
rect 583520 364784 584800 364896
rect 583520 363602 584800 363714
rect 2200 335050 18500 335250
rect 557250 362532 583550 362600
rect 557250 362420 584800 362532
rect 557250 362300 583550 362420
rect 557250 317100 560000 362300
rect 583520 361238 584800 361350
rect 583520 360056 584800 360168
rect 583520 358874 584800 358986
rect 583520 319562 584800 319674
rect 583520 318380 584800 318492
rect 483600 315100 560000 317100
rect 577700 317310 583650 317350
rect 577700 317198 584800 317310
rect 577700 317150 583650 317198
rect 577700 309100 579750 317150
rect 583520 316016 584800 316128
rect 583520 314834 584800 314946
rect 583520 313652 584800 313764
rect 483850 307950 579750 309100
rect 483850 307100 579550 307950
rect 1200 290800 3200 290850
rect 1200 290700 2950 290800
rect 3100 290700 3200 290800
rect 1200 290650 3200 290700
rect 583520 275140 584800 275252
rect 565450 274070 583550 274100
rect 565450 274050 584800 274070
rect 565450 273950 565500 274050
rect 565900 273958 584800 274050
rect 565900 273950 583550 273958
rect 565450 273900 583550 273950
rect 583520 272776 584800 272888
rect 583520 271594 584800 271706
rect 583520 270412 584800 270524
rect 583520 269230 584800 269342
rect 1200 248950 1850 249000
rect 1200 248850 1600 248950
rect 1750 248850 1850 248950
rect 1200 248800 1850 248850
rect 483450 233900 562500 235450
rect 582340 235230 584800 240030
rect 483550 228900 550950 230450
rect 1650 121400 1950 121450
rect 1400 121350 1950 121400
rect 1400 121250 1750 121350
rect 1900 121250 1950 121350
rect 1400 121200 1950 121250
rect 1650 121150 1950 121200
rect 1400 78100 2200 78150
rect 1400 78000 2000 78100
rect 2150 78000 2200 78100
rect 1400 77950 2200 78000
rect 549300 48250 550950 228900
rect 560950 92900 562500 233900
rect 582340 225230 584800 230030
rect 582340 191430 584800 196230
rect 582340 181430 584800 186230
rect 582340 146830 584800 151630
rect 582340 136830 584800 141630
rect 583520 95118 584800 95230
rect 583520 93936 584800 94048
rect 560950 92866 583600 92900
rect 560950 92754 584800 92866
rect 560950 92700 583600 92754
rect 583520 91572 584800 91684
rect 583520 50460 584800 50572
rect 583520 49278 584800 49390
rect 549300 48208 583550 48250
rect 549300 48096 584800 48208
rect 549300 48050 583550 48096
rect 583520 46914 584800 47026
rect 1400 34900 3350 34950
rect 1400 34800 3150 34900
rect 3300 34800 3350 34900
rect 1400 34750 3350 34800
<< via3 >>
rect 43280 689180 43860 690460
rect 45800 689180 46380 690460
rect 54174 688398 55256 688712
rect 57600 685400 58600 685600
rect 54202 682364 55256 682700
rect 5476 641552 8888 648570
rect 2434 557958 7216 563676
rect 263000 615000 263600 615800
rect 260800 613400 261400 614200
rect 302240 601140 302360 601240
rect 301820 597620 301980 597720
rect 333600 624000 334200 624800
rect 532800 624000 533600 624800
rect 307600 567000 307800 567200
rect 307600 566500 307800 566700
rect 2950 290700 3100 290800
rect 1600 248850 1750 248950
rect 1750 121250 1900 121350
rect 2000 78000 2150 78100
rect 3150 34800 3300 34900
<< metal4 >>
rect 165594 702300 170594 704800
rect 175894 702300 180894 704800
rect 217294 702300 222294 704800
rect 227594 702300 232594 704800
rect 318994 702300 323994 704800
rect 329294 702300 334294 704800
rect 43240 690460 44460 690500
rect 43240 689180 43280 690460
rect 43860 689180 44460 690460
rect 43240 689140 44460 689180
rect 44040 688220 44460 689140
rect 44720 690460 46460 690500
rect 44720 689180 45800 690460
rect 46380 689180 46460 690460
rect 44720 689140 46460 689180
rect 44720 688220 45140 689140
rect 54104 688712 55292 688744
rect 54104 688398 54174 688712
rect 55256 688398 55292 688712
rect 54104 682700 55292 688398
rect 54104 682364 54202 682700
rect 55256 682364 55292 682700
rect 47164 677302 47770 679332
rect 54104 677302 55292 682364
rect 47164 676830 55292 677302
rect 5062 648570 9348 648812
rect 5062 641552 5476 648570
rect 8888 641552 9348 648570
rect 5062 641230 9348 641552
rect 1636 563676 8000 564262
rect 1636 557958 2434 563676
rect 7216 557958 8000 563676
rect 1636 557296 8000 557958
rect 54104 563998 55292 676830
rect 57400 685600 58800 685800
rect 57400 685400 57600 685600
rect 58600 685400 58800 685600
rect 57400 614200 58800 685400
rect 177000 615800 180000 702300
rect 177000 615000 177200 615800
rect 179800 615000 180000 615800
rect 177000 614800 180000 615000
rect 232000 646000 237000 647000
rect 232000 643000 233000 646000
rect 236000 643000 237000 646000
rect 57400 613400 57600 614200
rect 58600 613400 58800 614200
rect 57400 613200 58800 613400
rect 232000 587400 237000 643000
rect 333599 624800 334201 624801
rect 333599 624000 333600 624800
rect 334200 624000 334201 624800
rect 333599 623999 334201 624000
rect 532799 624800 533601 624801
rect 532799 624000 532800 624800
rect 533600 624000 533601 624800
rect 532799 623999 533601 624000
rect 262999 615800 263601 615801
rect 262999 615000 263000 615800
rect 263600 615000 263601 615800
rect 262999 614999 263601 615000
rect 260799 614200 261401 614201
rect 260799 613400 260800 614200
rect 261400 613400 261401 614200
rect 260799 613399 261401 613400
rect 302200 601240 302400 601300
rect 302200 601140 302240 601240
rect 302360 601140 302400 601240
rect 301800 597720 302000 598000
rect 301800 597620 301820 597720
rect 301980 597620 302000 597720
rect 232000 586600 232800 587400
rect 236200 586600 240000 587400
rect 232000 586000 240000 586600
rect 54104 557596 54250 563998
rect 55084 557596 55292 563998
rect 238000 580300 239700 580800
rect 238000 562000 243000 580300
rect 238000 559000 239000 562000
rect 242000 559000 243000 562000
rect 238000 558000 243000 559000
rect 286000 562000 291000 580200
rect 301800 566700 302000 597620
rect 302200 567200 302400 601140
rect 307599 567200 307801 567201
rect 302200 567000 307600 567200
rect 307800 567000 307801 567200
rect 307599 566999 307801 567000
rect 307599 566700 307801 566701
rect 301800 566500 307600 566700
rect 307800 566500 307801 566700
rect 307599 566499 307801 566500
rect 286000 559000 287000 562000
rect 290000 559000 291000 562000
rect 298800 560200 306000 560400
rect 298800 559400 299000 560200
rect 299600 559400 306000 560200
rect 298800 559200 306000 559400
rect 286000 558000 291000 559000
rect 329200 558800 331200 560600
rect 329200 557800 329400 558800
rect 331000 557800 331200 558800
rect 329200 557600 331200 557800
rect 54104 557312 55292 557596
rect 2900 290800 96960 290950
rect 2900 290700 2950 290800
rect 3100 290700 96960 290800
rect 2900 290550 96960 290700
rect 1550 248950 37760 249100
rect 1550 248850 1600 248950
rect 1750 248850 37760 248950
rect 1550 248700 37760 248850
rect 37440 208960 37760 248700
rect 96640 218240 96960 290550
rect 37440 208920 87360 208960
rect 37440 208680 87080 208920
rect 87320 208680 87360 208920
rect 37440 208640 87360 208680
rect 37440 180120 89280 180160
rect 37440 179880 89000 180120
rect 89240 179880 89280 180120
rect 37440 179840 89280 179880
rect 37440 121450 37760 179840
rect 1700 121350 37760 121450
rect 1700 121250 1750 121350
rect 1900 121250 37760 121350
rect 1700 121150 37760 121250
rect 43520 158360 91840 158400
rect 43520 158120 91560 158360
rect 91800 158120 91840 158360
rect 43520 158080 91840 158120
rect 43520 78250 43840 158080
rect 1950 78100 43840 78250
rect 1950 78000 2000 78100
rect 2150 78000 43840 78100
rect 1950 77850 43840 78000
rect 48640 145880 94400 145920
rect 48640 145640 94120 145880
rect 94360 145640 94400 145880
rect 48640 145600 94400 145640
rect 48640 35050 48960 145600
rect 3100 34900 48960 35050
rect 3100 34800 3150 34900
rect 3300 34800 48960 34900
rect 3100 34650 48960 34800
<< via4 >>
rect 5476 641552 8888 648570
rect 2434 557958 7216 563676
rect 177200 615000 179800 615800
rect 233000 643000 236000 646000
rect 57600 613400 58600 614200
rect 333600 624000 334200 624800
rect 532800 624000 533600 624800
rect 263000 615000 263600 615800
rect 260800 613400 261400 614200
rect 232800 586600 236200 587400
rect 54250 557596 55084 563998
rect 239000 559000 242000 562000
rect 287000 559000 290000 562000
rect 299000 559400 299600 560200
rect 329400 557800 331000 558800
rect 87080 208680 87320 208920
rect 89000 179880 89240 180120
rect 91560 158120 91800 158360
rect 94120 145640 94360 145880
<< metal5 >>
rect 165594 702300 170594 704800
rect 175894 702300 180894 704800
rect 217294 702300 222294 704800
rect 227594 702300 232594 704800
rect 318994 702300 323994 704800
rect 329294 702300 334294 704800
rect 5062 648808 8864 648812
rect 42374 648808 42798 683446
rect 49922 648808 50564 683720
rect 5062 648570 305000 648808
rect 5062 641552 5476 648570
rect 8888 646000 305000 648570
rect 8888 643000 233000 646000
rect 236000 643000 305000 646000
rect 8888 641552 305000 643000
rect 5062 641230 305000 641552
rect 177000 615800 263800 616000
rect 177000 615000 177200 615800
rect 179800 615000 263000 615800
rect 263600 615000 263800 615800
rect 177000 614800 263800 615000
rect 57400 614200 261600 614400
rect 57400 613400 57600 614200
rect 58600 613400 260800 614200
rect 261400 613400 261600 614200
rect 57400 613200 261600 613400
rect 232600 587400 240000 587600
rect 232600 586600 232800 587400
rect 236200 586600 240000 587400
rect 232600 586400 240000 586600
rect 302800 565800 304200 641230
rect 333576 624800 334224 624824
rect 532776 624800 533624 624824
rect 333576 624000 333600 624800
rect 334200 624000 532800 624800
rect 533600 624000 533624 624800
rect 333576 623976 334224 624000
rect 532776 623976 533624 624000
rect 1636 563998 300000 564262
rect 1636 563676 54250 563998
rect 1636 557958 2434 563676
rect 7216 557958 54250 563676
rect 1636 557596 54250 557958
rect 55084 562000 300000 563998
rect 55084 559000 239000 562000
rect 242000 559000 287000 562000
rect 290000 560200 300000 562000
rect 290000 559400 299000 560200
rect 299600 559400 300000 560200
rect 290000 559296 300000 559400
rect 290000 559000 334000 559296
rect 55084 558800 334000 559000
rect 55084 557800 329400 558800
rect 331000 557800 334000 558800
rect 55084 557596 334000 557800
rect 1636 557296 334000 557596
<< comment >>
rect -100 704000 584100 704100
rect -100 0 0 704000
rect 584000 0 584100 704000
rect -100 -100 584100 0
use VCO-assembly  VCO-assembly_0
timestamp 1672466169
transform -1 0 60892 0 1 678180
box 6815 -326 25740 10562
use cmos_imager_rc_top  cmos_imager_rc_top_0
timestamp 1672454300
transform 1 0 305500 0 1 621000
box -1500 -61000 25600 28600
use current_ref  current_ref_0
timestamp 1672499013
transform 1 0 241000 0 1 581400
box -1400 -1400 52800 29800
use diode  diode_0
timestamp 1672465007
transform 1 0 570900 0 1 691340
box -200 -100 1210 796
use inductor_4  inductor_4_0
timestamp 1672460674
transform -1 0 97920 0 1 200960
box -17920 -62080 19840 35200
<< labels >>
flabel metal3 s 583520 269230 584800 269342 0 FreeSans 1120 0 0 0 gpio_analog[0]
port 0 nsew signal bidirectional
flabel metal3 s 583520 313652 584800 313764 0 FreeSans 1120 0 0 0 gpio_analog[1]
port 9 nsew signal bidirectional
flabel metal3 s 583520 358874 584800 358986 0 FreeSans 1120 0 0 0 gpio_analog[2]
port 10 nsew signal bidirectional
flabel metal3 s 583520 405296 584800 405408 0 FreeSans 1120 0 0 0 gpio_analog[3]
port 11 nsew signal bidirectional
flabel metal3 s 583520 449718 584800 449830 0 FreeSans 1120 0 0 0 gpio_analog[4]
port 12 nsew signal bidirectional
flabel metal3 s 583520 494140 584800 494252 0 FreeSans 1120 0 0 0 gpio_analog[5]
port 13 nsew signal bidirectional
flabel metal3 s 583520 583562 584800 583674 0 FreeSans 1120 0 0 0 gpio_analog[6]
port 14 nsew signal bidirectional
flabel metal3 s 583520 270412 584800 270524 0 FreeSans 1120 0 0 0 gpio_noesd[0]
port 18 nsew signal bidirectional
flabel metal3 s 583520 314834 584800 314946 0 FreeSans 1120 0 0 0 gpio_noesd[1]
port 27 nsew signal bidirectional
flabel metal3 s 583520 360056 584800 360168 0 FreeSans 1120 0 0 0 gpio_noesd[2]
port 28 nsew signal bidirectional
flabel metal3 s 583520 406478 584800 406590 0 FreeSans 1120 0 0 0 gpio_noesd[3]
port 29 nsew signal bidirectional
flabel metal3 s 583520 450900 584800 451012 0 FreeSans 1120 0 0 0 gpio_noesd[4]
port 30 nsew signal bidirectional
flabel metal3 s 583520 495322 584800 495434 0 FreeSans 1120 0 0 0 gpio_noesd[5]
port 31 nsew signal bidirectional
flabel metal3 s 583520 584744 584800 584856 0 FreeSans 1120 0 0 0 gpio_noesd[6]
port 32 nsew signal bidirectional
flabel metal3 s 582300 677984 584800 682984 0 FreeSans 1120 0 0 0 io_analog[0]
port 36 nsew signal bidirectional
flabel metal3 s 566594 702300 571594 704800 0 FreeSans 1920 180 0 0 io_analog[1]
port 38 nsew signal bidirectional
flabel metal3 s 465394 702300 470394 704800 0 FreeSans 1920 180 0 0 io_analog[2]
port 39 nsew signal bidirectional
flabel metal3 s 413394 702300 418394 704800 0 FreeSans 1920 180 0 0 io_analog[3]
port 40 nsew signal bidirectional
flabel metal3 s 329294 702300 334294 704800 0 FreeSans 1920 180 0 0 io_analog[4]
port 41 nsew signal bidirectional
flabel metal4 s 329294 702300 334294 704800 0 FreeSans 1920 180 0 0 io_analog[4]
port 41 nsew signal bidirectional
flabel metal5 s 329294 702300 334294 704800 0 FreeSans 1920 180 0 0 io_analog[4]
port 41 nsew signal bidirectional
flabel metal3 s 227594 702300 232594 704800 0 FreeSans 1920 180 0 0 io_analog[5]
port 42 nsew signal bidirectional
flabel metal4 s 227594 702300 232594 704800 0 FreeSans 1920 180 0 0 io_analog[5]
port 42 nsew signal bidirectional
flabel metal5 s 227594 702300 232594 704800 0 FreeSans 1920 180 0 0 io_analog[5]
port 42 nsew signal bidirectional
flabel metal3 s 175894 702300 180894 704800 0 FreeSans 1920 180 0 0 io_analog[6]
port 43 nsew signal bidirectional
flabel metal4 s 175894 702300 180894 704800 0 FreeSans 1920 180 0 0 io_analog[6]
port 43 nsew signal bidirectional
flabel metal5 s 175894 702300 180894 704800 0 FreeSans 1920 180 0 0 io_analog[6]
port 43 nsew signal bidirectional
flabel metal3 s 120194 702300 125194 704800 0 FreeSans 1920 180 0 0 io_analog[7]
port 44 nsew signal bidirectional
flabel metal3 s 318994 702300 323994 704800 0 FreeSans 1920 180 0 0 io_analog[4]
port 47 nsew signal bidirectional
flabel metal4 s 318994 702300 323994 704800 0 FreeSans 1920 180 0 0 io_analog[4]
port 47 nsew signal bidirectional
flabel metal5 s 318994 702300 323994 704800 0 FreeSans 1920 180 0 0 io_analog[4]
port 47 nsew signal bidirectional
flabel metal3 s 217294 702300 222294 704800 0 FreeSans 1920 180 0 0 io_analog[5]
port 48 nsew signal bidirectional
flabel metal4 s 217294 702300 222294 704800 0 FreeSans 1920 180 0 0 io_analog[5]
port 48 nsew signal bidirectional
flabel metal5 s 217294 702300 222294 704800 0 FreeSans 1920 180 0 0 io_analog[5]
port 48 nsew signal bidirectional
flabel metal3 s 165594 702300 170594 704800 0 FreeSans 1920 180 0 0 io_analog[6]
port 49 nsew signal bidirectional
flabel metal4 s 165594 702300 170594 704800 0 FreeSans 1920 180 0 0 io_analog[6]
port 49 nsew signal bidirectional
flabel metal5 s 165594 702300 170594 704800 0 FreeSans 1920 180 0 0 io_analog[6]
port 49 nsew signal bidirectional
flabel metal3 s 326794 702300 328994 704800 0 FreeSans 1920 180 0 0 io_clamp_high[0]
port 50 nsew signal bidirectional
flabel metal3 s 225094 702300 227294 704800 0 FreeSans 1920 180 0 0 io_clamp_high[1]
port 51 nsew signal bidirectional
flabel metal3 s 173394 702300 175594 704800 0 FreeSans 1920 180 0 0 io_clamp_high[2]
port 52 nsew signal bidirectional
flabel metal3 s 324294 702300 326494 704800 0 FreeSans 1920 180 0 0 io_clamp_low[0]
port 53 nsew signal bidirectional
flabel metal3 s 222594 702300 224794 704800 0 FreeSans 1920 180 0 0 io_clamp_low[1]
port 54 nsew signal bidirectional
flabel metal3 s 170894 702300 173094 704800 0 FreeSans 1920 180 0 0 io_clamp_low[2]
port 55 nsew signal bidirectional
flabel metal3 s 583520 408842 584800 408954 0 FreeSans 1120 0 0 0 io_in[10]
port 57 nsew signal input
flabel metal3 s 583520 453264 584800 453376 0 FreeSans 1120 0 0 0 io_in[11]
port 58 nsew signal input
flabel metal3 s 583520 497686 584800 497798 0 FreeSans 1120 0 0 0 io_in[12]
port 59 nsew signal input
flabel metal3 s 583520 587108 584800 587220 0 FreeSans 1120 0 0 0 io_in[13]
port 60 nsew signal input
flabel metal3 s 583520 48096 584800 48208 0 FreeSans 1120 0 0 0 io_in[5]
port 78 nsew signal input
flabel metal3 s 583520 92754 584800 92866 0 FreeSans 1120 0 0 0 io_in[6]
port 79 nsew signal input
flabel metal3 s 583520 272776 584800 272888 0 FreeSans 1120 0 0 0 io_in[7]
port 80 nsew signal input
flabel metal3 s 583520 317198 584800 317310 0 FreeSans 1120 0 0 0 io_in[8]
port 81 nsew signal input
flabel metal3 s 583520 362420 584800 362532 0 FreeSans 1120 0 0 0 io_in[9]
port 82 nsew signal input
flabel metal3 s 583520 407660 584800 407772 0 FreeSans 1120 0 0 0 io_in_3v3[10]
port 84 nsew signal input
flabel metal3 s 583520 452082 584800 452194 0 FreeSans 1120 0 0 0 io_in_3v3[11]
port 85 nsew signal input
flabel metal3 s 583520 496504 584800 496616 0 FreeSans 1120 0 0 0 io_in_3v3[12]
port 86 nsew signal input
flabel metal3 s 583520 585926 584800 586038 0 FreeSans 1120 0 0 0 io_in_3v3[13]
port 87 nsew signal input
flabel metal3 s 583520 46914 584800 47026 0 FreeSans 1120 0 0 0 io_in_3v3[5]
port 105 nsew signal input
flabel metal3 s 583520 91572 584800 91684 0 FreeSans 1120 0 0 0 io_in_3v3[6]
port 106 nsew signal input
flabel metal3 s 583520 271594 584800 271706 0 FreeSans 1120 0 0 0 io_in_3v3[7]
port 107 nsew signal input
flabel metal3 s 583520 316016 584800 316128 0 FreeSans 1120 0 0 0 io_in_3v3[8]
port 108 nsew signal input
flabel metal3 s 583520 361238 584800 361350 0 FreeSans 1120 0 0 0 io_in_3v3[9]
port 109 nsew signal input
flabel metal3 s 583520 411206 584800 411318 0 FreeSans 1120 0 0 0 io_oeb[10]
port 111 nsew signal tristate
flabel metal3 s 583520 455628 584800 455740 0 FreeSans 1120 0 0 0 io_oeb[11]
port 112 nsew signal tristate
flabel metal3 s 583520 500050 584800 500162 0 FreeSans 1120 0 0 0 io_oeb[12]
port 113 nsew signal tristate
flabel metal3 s 583520 589472 584800 589584 0 FreeSans 1120 0 0 0 io_oeb[13]
port 114 nsew signal tristate
flabel metal3 s 583520 50460 584800 50572 0 FreeSans 1120 0 0 0 io_oeb[5]
port 132 nsew signal tristate
flabel metal3 s 583520 95118 584800 95230 0 FreeSans 1120 0 0 0 io_oeb[6]
port 133 nsew signal tristate
flabel metal3 s 583520 275140 584800 275252 0 FreeSans 1120 0 0 0 io_oeb[7]
port 134 nsew signal tristate
flabel metal3 s 583520 319562 584800 319674 0 FreeSans 1120 0 0 0 io_oeb[8]
port 135 nsew signal tristate
flabel metal3 s 583520 364784 584800 364896 0 FreeSans 1120 0 0 0 io_oeb[9]
port 136 nsew signal tristate
flabel metal3 s 583520 410024 584800 410136 0 FreeSans 1120 0 0 0 io_out[10]
port 138 nsew signal tristate
flabel metal3 s 583520 454446 584800 454558 0 FreeSans 1120 0 0 0 io_out[11]
port 139 nsew signal tristate
flabel metal3 s 583520 498868 584800 498980 0 FreeSans 1120 0 0 0 io_out[12]
port 140 nsew signal tristate
flabel metal3 s 583520 588290 584800 588402 0 FreeSans 1120 0 0 0 io_out[13]
port 141 nsew signal tristate
flabel metal3 s 583520 49278 584800 49390 0 FreeSans 1120 0 0 0 io_out[5]
port 159 nsew signal tristate
flabel metal3 s 583520 93936 584800 94048 0 FreeSans 1120 0 0 0 io_out[6]
port 160 nsew signal tristate
flabel metal3 s 583520 273958 584800 274070 0 FreeSans 1120 0 0 0 io_out[7]
port 161 nsew signal tristate
flabel metal3 s 583520 318380 584800 318492 0 FreeSans 1120 0 0 0 io_out[8]
port 162 nsew signal tristate
flabel metal3 s 583520 363602 584800 363714 0 FreeSans 1120 0 0 0 io_out[9]
port 163 nsew signal tristate
flabel metal3 s 582340 639784 584800 644584 0 FreeSans 1120 0 0 0 vccd1
port 552 nsew signal bidirectional
flabel metal3 s 582340 629784 584800 634584 0 FreeSans 1120 0 0 0 vccd1
port 553 nsew signal bidirectional
flabel metal3 s 582340 540562 584800 545362 0 FreeSans 1120 0 0 0 vdda1
port 556 nsew signal bidirectional
flabel metal3 s 582340 550562 584800 555362 0 FreeSans 1120 0 0 0 vdda1
port 557 nsew signal bidirectional
flabel metal3 s 582340 235230 584800 240030 0 FreeSans 1120 0 0 0 vdda1
port 558 nsew signal bidirectional
flabel metal3 s 582340 225230 584800 230030 0 FreeSans 1120 0 0 0 vdda1
port 559 nsew signal bidirectional
flabel metal3 s 520594 702340 525394 704800 0 FreeSans 1920 180 0 0 vssa1
port 562 nsew signal bidirectional
flabel metal3 s 510594 702340 515394 704800 0 FreeSans 1920 180 0 0 vssa1
port 563 nsew signal bidirectional
flabel metal3 s 582340 146830 584800 151630 0 FreeSans 1120 0 0 0 vssa1
port 564 nsew signal bidirectional
flabel metal3 s 582340 136830 584800 141630 0 FreeSans 1120 0 0 0 vssa1
port 565 nsew signal bidirectional
flabel metal3 s 582340 191430 584800 196230 0 FreeSans 1120 0 0 0 vssd1
port 568 nsew signal bidirectional
flabel metal3 s 582340 181430 584800 186230 0 FreeSans 1120 0 0 0 vssd1
port 569 nsew signal bidirectional
flabel space 52726 685400 56918 685476 3 FreeSans 1600 0 0 0 BIAS
flabel space 474800 417000 512000 430200 0 FreeSans 80000 0 0 0 sh_clk
flabel space 471600 459900 512600 466900 0 FreeSans 80000 0 0 0 B
flabel space 472000 502400 513000 509400 0 FreeSans 80000 0 0 0 A
flabel space 90700 617200 104500 622000 0 FreeSans 80000 0 0 0 I=40uA
flabel space 126300 688300 140100 693100 0 FreeSans 80000 0 0 0 Vbg
flabel space 248000 657000 265000 663000 0 FreeSans 64000 0 0 0 RC_Imager_Out
flabel space 503000 627400 512800 630000 0 FreeSans 64000 0 0 0 rst_b_clk
<< properties >>
string FIXED_BBOX 0 0 584000 704000
<< end >>
