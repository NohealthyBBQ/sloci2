magic
tech sky130A
magscale 1 2
timestamp 1672435296
<< locali >>
rect 11660 5680 16200 5740
rect 11660 5420 16200 5490
rect 11660 5240 16210 5290
rect 11660 4990 16210 5040
rect 11720 4500 13100 4660
rect 14760 4500 16140 4660
rect 11720 4220 13100 4380
rect 14760 4220 16140 4380
rect 11660 3840 16210 3890
rect 11660 3590 16210 3640
rect 11670 3390 16220 3440
rect 11660 3140 16210 3190
<< metal1 >>
rect 11790 2650 13030 2710
rect 12390 2340 12440 2650
rect 11790 2290 13030 2340
rect 38410 -320 38420 -100
rect 38800 -320 38810 -100
rect 27630 -840 27640 -620
rect 28000 -840 28010 -620
<< via1 >>
rect 38420 -320 38800 -100
rect 27640 -840 28000 -620
<< metal2 >>
rect 7300 3000 11400 3200
rect 1700 1860 1800 1870
rect 1700 1750 1800 1760
rect 2160 1860 2280 1880
rect 2160 1760 2170 1860
rect 2260 1760 2280 1860
rect 2160 1680 2280 1760
rect 2160 1580 2880 1680
rect 38400 -100 38820 -80
rect 38400 -320 38420 -100
rect 38800 -320 38820 -100
rect 38400 -500 38820 -320
rect 27640 -620 38820 -500
rect 28000 -840 38820 -620
rect 27640 -960 38820 -840
<< via2 >>
rect 1700 1760 1800 1860
rect 2170 1760 2260 1860
<< metal3 >>
rect 1690 1860 2270 1870
rect 1690 1760 1700 1860
rect 1800 1760 2170 1860
rect 2260 1760 2270 1860
rect 1690 1750 2270 1760
use XM_Rref  XM_Rref_0
timestamp 1662826901
transform 0 1 18173 1 0 1417
box -1417 -1173 5029 21223
use XM_current_gate_with_dummy  XM_current_gate_with_dummy_0
timestamp 1662842659
transform 1 0 11600 0 1 3924
box 0 -924 4660 1954
use XM_output_mirr_combined_with_dummy  XM_output_mirr_combined_with_dummy_0
timestamp 1662903677
transform 1 0 16600 0 1 14200
box -17600 -7400 35500 15000
use opamp_realcomp3_usefinger  opamp_realcomp3_usefinger_0
timestamp 1662836520
transform 1 0 4380 0 1 -594
box -5380 594 6776 6403
use sky130_fd_pr__nfet_01v8_lvt_E2U6GT  sky130_fd_pr__nfet_01v8_lvt_E2U6GT_0
timestamp 1672431769
transform 1 0 12196 0 1 1359
box -596 -679 596 679
use sky130_fd_pr__nfet_01v8_lvt_H8V8HY  sky130_fd_pr__nfet_01v8_lvt_H8V8HY_0
timestamp 1672431769
transform 1 0 13096 0 1 859
box -396 -1179 396 1179
use sky130_fd_pr__pfet_01v8_lvt_MUVN4U  sky130_fd_pr__pfet_01v8_lvt_MUVN4U_0
timestamp 1672432293
transform 1 0 12412 0 1 2626
box -812 -466 812 466
use sky130_fd_pr__res_high_po_1p41_EL7NMZ  sky130_fd_pr__res_high_po_1p41_EL7NMZ_0
timestamp 1672432498
transform 0 -1 22598 1 0 -733
box -307 -5598 307 5598
use sky130_fd_pr__res_high_po_1p41_G3LFBQ  sky130_fd_pr__res_high_po_1p41_G3LFBQ_0
timestamp 1672432498
transform 0 1 27998 -1 0 -213
box -307 -10998 307 10998
<< labels >>
flabel space 13210 4940 13250 5000 0 FreeSans 960 0 0 0 C
flabel space 14620 4940 14660 5000 0 FreeSans 960 0 0 0 C
flabel space 13200 3850 13240 3910 0 FreeSans 960 0 0 0 C
flabel space 14620 3870 14660 3930 0 FreeSans 960 0 0 0 C
<< end >>
