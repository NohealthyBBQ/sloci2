magic
tech sky130A
magscale 1 2
timestamp 1662720466
<< nwell >>
rect -812 -466 812 466
<< pmoslvt >>
rect -616 118 -416 318
rect -358 118 -158 318
rect -100 118 100 318
rect 158 118 358 318
rect 416 118 616 318
rect -616 -247 -416 -47
rect -358 -247 -158 -47
rect -100 -247 100 -47
rect 158 -247 358 -47
rect 416 -247 616 -47
<< pdiff >>
rect -674 306 -616 318
rect -674 130 -662 306
rect -628 130 -616 306
rect -674 118 -616 130
rect -416 306 -358 318
rect -416 130 -404 306
rect -370 130 -358 306
rect -416 118 -358 130
rect -158 306 -100 318
rect -158 130 -146 306
rect -112 130 -100 306
rect -158 118 -100 130
rect 100 306 158 318
rect 100 130 112 306
rect 146 130 158 306
rect 100 118 158 130
rect 358 306 416 318
rect 358 130 370 306
rect 404 130 416 306
rect 358 118 416 130
rect 616 306 674 318
rect 616 130 628 306
rect 662 130 674 306
rect 616 118 674 130
rect -674 -59 -616 -47
rect -674 -235 -662 -59
rect -628 -235 -616 -59
rect -674 -247 -616 -235
rect -416 -59 -358 -47
rect -416 -235 -404 -59
rect -370 -235 -358 -59
rect -416 -247 -358 -235
rect -158 -59 -100 -47
rect -158 -235 -146 -59
rect -112 -235 -100 -59
rect -158 -247 -100 -235
rect 100 -59 158 -47
rect 100 -235 112 -59
rect 146 -235 158 -59
rect 100 -247 158 -235
rect 358 -59 416 -47
rect 358 -235 370 -59
rect 404 -235 416 -59
rect 358 -247 416 -235
rect 616 -59 674 -47
rect 616 -235 628 -59
rect 662 -235 674 -59
rect 616 -247 674 -235
<< pdiffc >>
rect -662 130 -628 306
rect -404 130 -370 306
rect -146 130 -112 306
rect 112 130 146 306
rect 370 130 404 306
rect 628 130 662 306
rect -662 -235 -628 -59
rect -404 -235 -370 -59
rect -146 -235 -112 -59
rect 112 -235 146 -59
rect 370 -235 404 -59
rect 628 -235 662 -59
<< nsubdiff >>
rect -776 396 -680 430
rect 680 396 776 430
rect -776 334 -742 396
rect 742 334 776 396
rect -776 -396 -742 -334
rect 742 -396 776 -334
rect -776 -430 -680 -396
rect 680 -430 776 -396
<< nsubdiffcont >>
rect -680 396 680 430
rect -776 -334 -742 334
rect 742 -334 776 334
rect -680 -430 680 -396
<< poly >>
rect -616 318 -416 344
rect -358 318 -158 344
rect -100 318 100 344
rect 158 318 358 344
rect 416 318 616 344
rect -616 71 -416 118
rect -616 37 -600 71
rect -432 37 -416 71
rect -616 21 -416 37
rect -358 71 -158 118
rect -358 37 -342 71
rect -174 37 -158 71
rect -358 21 -158 37
rect -100 71 100 118
rect -100 37 -84 71
rect 84 37 100 71
rect -100 21 100 37
rect 158 71 358 118
rect 158 37 174 71
rect 342 37 358 71
rect 158 21 358 37
rect 416 71 616 118
rect 416 37 432 71
rect 600 37 616 71
rect 416 21 616 37
rect -616 -47 -416 -21
rect -358 -47 -158 -21
rect -100 -47 100 -21
rect 158 -47 358 -21
rect 416 -47 616 -21
rect -616 -294 -416 -247
rect -616 -328 -600 -294
rect -432 -328 -416 -294
rect -616 -344 -416 -328
rect -358 -294 -158 -247
rect -358 -328 -342 -294
rect -174 -328 -158 -294
rect -358 -344 -158 -328
rect -100 -294 100 -247
rect -100 -328 -84 -294
rect 84 -328 100 -294
rect -100 -344 100 -328
rect 158 -294 358 -247
rect 158 -328 174 -294
rect 342 -328 358 -294
rect 158 -344 358 -328
rect 416 -294 616 -247
rect 416 -328 432 -294
rect 600 -328 616 -294
rect 416 -344 616 -328
<< polycont >>
rect -600 37 -432 71
rect -342 37 -174 71
rect -84 37 84 71
rect 174 37 342 71
rect 432 37 600 71
rect -600 -328 -432 -294
rect -342 -328 -174 -294
rect -84 -328 84 -294
rect 174 -328 342 -294
rect 432 -328 600 -294
<< locali >>
rect -776 396 -680 430
rect 680 396 776 430
rect -776 334 -742 396
rect 742 334 776 396
rect -662 306 -628 322
rect -662 114 -628 130
rect -404 306 -370 322
rect -404 114 -370 130
rect -146 306 -112 322
rect -146 114 -112 130
rect 112 306 146 322
rect 112 114 146 130
rect 370 306 404 322
rect 370 114 404 130
rect 628 306 662 322
rect 628 114 662 130
rect -616 37 -600 71
rect -432 37 -416 71
rect -358 37 -342 71
rect -174 37 -158 71
rect -100 37 -84 71
rect 84 37 100 71
rect 158 37 174 71
rect 342 37 358 71
rect 416 37 432 71
rect 600 37 616 71
rect -662 -59 -628 -43
rect -662 -251 -628 -235
rect -404 -59 -370 -43
rect -404 -251 -370 -235
rect -146 -59 -112 -43
rect -146 -251 -112 -235
rect 112 -59 146 -43
rect 112 -251 146 -235
rect 370 -59 404 -43
rect 370 -251 404 -235
rect 628 -59 662 -43
rect 628 -251 662 -235
rect -616 -328 -600 -294
rect -432 -328 -416 -294
rect -358 -328 -342 -294
rect -174 -328 -158 -294
rect -100 -328 -84 -294
rect 84 -328 100 -294
rect 158 -328 174 -294
rect 342 -328 358 -294
rect 416 -328 432 -294
rect 600 -328 616 -294
rect -776 -396 -742 -334
rect 742 -396 776 -334
rect -776 -430 -680 -396
rect 680 -430 776 -396
<< viali >>
rect -662 130 -628 306
rect -404 130 -370 306
rect -146 130 -112 306
rect 112 130 146 306
rect 370 130 404 306
rect 628 130 662 306
rect -600 37 -432 71
rect -342 37 -174 71
rect -84 37 84 71
rect 174 37 342 71
rect 432 37 600 71
rect -662 -235 -628 -59
rect -404 -235 -370 -59
rect -146 -235 -112 -59
rect 112 -235 146 -59
rect 370 -235 404 -59
rect 628 -235 662 -59
rect -600 -328 -432 -294
rect -342 -328 -174 -294
rect -84 -328 84 -294
rect 174 -328 342 -294
rect 432 -328 600 -294
<< metal1 >>
rect -668 306 -622 318
rect -668 130 -662 306
rect -628 130 -622 306
rect -668 118 -622 130
rect -410 306 -364 318
rect -410 130 -404 306
rect -370 130 -364 306
rect -410 118 -364 130
rect -152 306 -106 318
rect -152 130 -146 306
rect -112 130 -106 306
rect -152 118 -106 130
rect 106 306 152 318
rect 106 130 112 306
rect 146 130 152 306
rect 106 118 152 130
rect 364 306 410 318
rect 364 130 370 306
rect 404 130 410 306
rect 364 118 410 130
rect 622 306 668 318
rect 622 130 628 306
rect 662 130 668 306
rect 622 118 668 130
rect -612 71 -420 77
rect -612 37 -600 71
rect -432 37 -420 71
rect -612 31 -420 37
rect -354 71 -162 77
rect -354 37 -342 71
rect -174 37 -162 71
rect -354 31 -162 37
rect -96 71 96 77
rect -96 37 -84 71
rect 84 37 96 71
rect -96 31 96 37
rect 162 71 354 77
rect 162 37 174 71
rect 342 37 354 71
rect 162 31 354 37
rect 420 71 612 77
rect 420 37 432 71
rect 600 37 612 71
rect 420 31 612 37
rect -668 -59 -622 -47
rect -668 -235 -662 -59
rect -628 -235 -622 -59
rect -668 -247 -622 -235
rect -410 -59 -364 -47
rect -410 -235 -404 -59
rect -370 -235 -364 -59
rect -410 -247 -364 -235
rect -152 -59 -106 -47
rect -152 -235 -146 -59
rect -112 -235 -106 -59
rect -152 -247 -106 -235
rect 106 -59 152 -47
rect 106 -235 112 -59
rect 146 -235 152 -59
rect 106 -247 152 -235
rect 364 -59 410 -47
rect 364 -235 370 -59
rect 404 -235 410 -59
rect 364 -247 410 -235
rect 622 -59 668 -47
rect 622 -235 628 -59
rect 662 -235 668 -59
rect 622 -247 668 -235
rect -612 -294 -420 -288
rect -612 -328 -600 -294
rect -432 -328 -420 -294
rect -612 -334 -420 -328
rect -354 -294 -162 -288
rect -354 -328 -342 -294
rect -174 -328 -162 -294
rect -354 -334 -162 -328
rect -96 -294 96 -288
rect -96 -328 -84 -294
rect 84 -328 96 -294
rect -96 -334 96 -328
rect 162 -294 354 -288
rect 162 -328 174 -294
rect 342 -328 354 -294
rect 162 -334 354 -328
rect 420 -294 612 -288
rect 420 -328 432 -294
rect 600 -328 612 -294
rect 420 -334 612 -328
<< properties >>
string FIXED_BBOX -759 -413 759 413
string gencell sky130_fd_pr__pfet_01v8_lvt
string library sky130
string parameters w 1 l 1 m 2 nf 5 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 0 botc 1 poverlap 0 doverlap 1 lmin 0.35 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
