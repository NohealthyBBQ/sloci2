magic
tech sky130A
magscale 1 2
timestamp 1672279567
<< metal3 >>
rect -3150 12522 3149 12550
rect -3150 6378 3065 12522
rect 3129 6378 3149 12522
rect -3150 6350 3149 6378
rect -3150 6222 3149 6250
rect -3150 78 3065 6222
rect 3129 78 3149 6222
rect -3150 50 3149 78
rect -3150 -78 3149 -50
rect -3150 -6222 3065 -78
rect 3129 -6222 3149 -78
rect -3150 -6250 3149 -6222
rect -3150 -6378 3149 -6350
rect -3150 -12522 3065 -6378
rect 3129 -12522 3149 -6378
rect -3150 -12550 3149 -12522
<< via3 >>
rect 3065 6378 3129 12522
rect 3065 78 3129 6222
rect 3065 -6222 3129 -78
rect 3065 -12522 3129 -6378
<< mimcap >>
rect -3050 12410 2950 12450
rect -3050 6490 -3010 12410
rect 2910 6490 2950 12410
rect -3050 6450 2950 6490
rect -3050 6110 2950 6150
rect -3050 190 -3010 6110
rect 2910 190 2950 6110
rect -3050 150 2950 190
rect -3050 -190 2950 -150
rect -3050 -6110 -3010 -190
rect 2910 -6110 2950 -190
rect -3050 -6150 2950 -6110
rect -3050 -6490 2950 -6450
rect -3050 -12410 -3010 -6490
rect 2910 -12410 2950 -6490
rect -3050 -12450 2950 -12410
<< mimcapcontact >>
rect -3010 6490 2910 12410
rect -3010 190 2910 6110
rect -3010 -6110 2910 -190
rect -3010 -12410 2910 -6490
<< metal4 >>
rect -102 12411 2 12600
rect 3018 12538 3122 12600
rect 3018 12522 3145 12538
rect -3011 12410 2911 12411
rect -3011 6490 -3010 12410
rect 2910 6490 2911 12410
rect -3011 6489 2911 6490
rect -102 6111 2 6489
rect 3018 6378 3065 12522
rect 3129 6378 3145 12522
rect 3018 6362 3145 6378
rect 3018 6238 3122 6362
rect 3018 6222 3145 6238
rect -3011 6110 2911 6111
rect -3011 190 -3010 6110
rect 2910 190 2911 6110
rect -3011 189 2911 190
rect -102 -189 2 189
rect 3018 78 3065 6222
rect 3129 78 3145 6222
rect 3018 62 3145 78
rect 3018 -62 3122 62
rect 3018 -78 3145 -62
rect -3011 -190 2911 -189
rect -3011 -6110 -3010 -190
rect 2910 -6110 2911 -190
rect -3011 -6111 2911 -6110
rect -102 -6489 2 -6111
rect 3018 -6222 3065 -78
rect 3129 -6222 3145 -78
rect 3018 -6238 3145 -6222
rect 3018 -6362 3122 -6238
rect 3018 -6378 3145 -6362
rect -3011 -6490 2911 -6489
rect -3011 -12410 -3010 -6490
rect 2910 -12410 2911 -6490
rect -3011 -12411 2911 -12410
rect -102 -12600 2 -12411
rect 3018 -12522 3065 -6378
rect 3129 -12522 3145 -6378
rect 3018 -12538 3145 -12522
rect 3018 -12600 3122 -12538
<< properties >>
string FIXED_BBOX -3150 6350 3050 12550
string gencell sky130_fd_pr__cap_mim_m3_1
string library sky130
string parameters w 30 l 30 val 1.822k carea 2.00 cperi 0.19 nx 1 ny 4 dummy 0 square 0 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 1 tconnect 1 ccov 100
<< end >>
