magic
tech sky130A
magscale 1 2
timestamp 1662765605
<< pwell >>
rect -1083 -1857 1083 1857
<< nmoslvt >>
rect -887 109 -487 1709
rect -429 109 -29 1709
rect 29 109 429 1709
rect 487 109 887 1709
rect -887 -1647 -487 -47
rect -429 -1647 -29 -47
rect 29 -1647 429 -47
rect 487 -1647 887 -47
<< ndiff >>
rect -945 1697 -887 1709
rect -945 121 -933 1697
rect -899 121 -887 1697
rect -945 109 -887 121
rect -487 1697 -429 1709
rect -487 121 -475 1697
rect -441 121 -429 1697
rect -487 109 -429 121
rect -29 1697 29 1709
rect -29 121 -17 1697
rect 17 121 29 1697
rect -29 109 29 121
rect 429 1697 487 1709
rect 429 121 441 1697
rect 475 121 487 1697
rect 429 109 487 121
rect 887 1697 945 1709
rect 887 121 899 1697
rect 933 121 945 1697
rect 887 109 945 121
rect -945 -59 -887 -47
rect -945 -1635 -933 -59
rect -899 -1635 -887 -59
rect -945 -1647 -887 -1635
rect -487 -59 -429 -47
rect -487 -1635 -475 -59
rect -441 -1635 -429 -59
rect -487 -1647 -429 -1635
rect -29 -59 29 -47
rect -29 -1635 -17 -59
rect 17 -1635 29 -59
rect -29 -1647 29 -1635
rect 429 -59 487 -47
rect 429 -1635 441 -59
rect 475 -1635 487 -59
rect 429 -1647 487 -1635
rect 887 -59 945 -47
rect 887 -1635 899 -59
rect 933 -1635 945 -59
rect 887 -1647 945 -1635
<< ndiffc >>
rect -933 121 -899 1697
rect -475 121 -441 1697
rect -17 121 17 1697
rect 441 121 475 1697
rect 899 121 933 1697
rect -933 -1635 -899 -59
rect -475 -1635 -441 -59
rect -17 -1635 17 -59
rect 441 -1635 475 -59
rect 899 -1635 933 -59
<< psubdiff >>
rect -1047 1787 -951 1821
rect 951 1787 1047 1821
rect -1047 -1787 -1013 1787
rect 1013 -1787 1047 1787
rect -1047 -1821 -951 -1787
rect 951 -1821 1047 -1787
<< psubdiffcont >>
rect -951 1787 951 1821
rect -951 -1821 951 -1787
<< poly >>
rect -887 1709 -487 1735
rect -429 1709 -29 1735
rect 29 1709 429 1735
rect 487 1709 887 1735
rect -887 71 -487 109
rect -887 37 -871 71
rect -503 37 -487 71
rect -887 21 -487 37
rect -429 71 -29 109
rect -429 37 -413 71
rect -45 37 -29 71
rect -429 21 -29 37
rect 29 71 429 109
rect 29 37 45 71
rect 413 37 429 71
rect 29 21 429 37
rect 487 71 887 109
rect 487 37 503 71
rect 871 37 887 71
rect 487 21 887 37
rect -887 -47 -487 -21
rect -429 -47 -29 -21
rect 29 -47 429 -21
rect 487 -47 887 -21
rect -887 -1685 -487 -1647
rect -887 -1719 -871 -1685
rect -503 -1719 -487 -1685
rect -887 -1735 -487 -1719
rect -429 -1685 -29 -1647
rect -429 -1719 -413 -1685
rect -45 -1719 -29 -1685
rect -429 -1735 -29 -1719
rect 29 -1685 429 -1647
rect 29 -1719 45 -1685
rect 413 -1719 429 -1685
rect 29 -1735 429 -1719
rect 487 -1685 887 -1647
rect 487 -1719 503 -1685
rect 871 -1719 887 -1685
rect 487 -1735 887 -1719
<< polycont >>
rect -871 37 -503 71
rect -413 37 -45 71
rect 45 37 413 71
rect 503 37 871 71
rect -871 -1719 -503 -1685
rect -413 -1719 -45 -1685
rect 45 -1719 413 -1685
rect 503 -1719 871 -1685
<< locali >>
rect -1047 1787 -951 1821
rect 951 1787 1047 1821
rect -1047 -1787 -1013 1787
rect -933 1697 -899 1713
rect -933 105 -899 121
rect -475 1697 -441 1713
rect -475 105 -441 121
rect -17 1697 17 1713
rect -17 105 17 121
rect 441 1697 475 1713
rect 441 105 475 121
rect 899 1697 933 1713
rect 899 105 933 121
rect -887 37 -871 71
rect -503 37 -487 71
rect -429 37 -413 71
rect -45 37 -29 71
rect 29 37 45 71
rect 413 37 429 71
rect 487 37 503 71
rect 871 37 887 71
rect -933 -59 -899 -43
rect -933 -1651 -899 -1635
rect -475 -59 -441 -43
rect -475 -1651 -441 -1635
rect -17 -59 17 -43
rect -17 -1651 17 -1635
rect 441 -59 475 -43
rect 441 -1651 475 -1635
rect 899 -59 933 -43
rect 899 -1651 933 -1635
rect -887 -1719 -871 -1685
rect -503 -1719 -487 -1685
rect -429 -1719 -413 -1685
rect -45 -1719 -29 -1685
rect 29 -1719 45 -1685
rect 413 -1719 429 -1685
rect 487 -1719 503 -1685
rect 871 -1719 887 -1685
rect 1013 -1787 1047 1787
rect -1047 -1821 -951 -1787
rect 951 -1821 1047 -1787
<< viali >>
rect -933 121 -899 1697
rect -475 121 -441 1697
rect -17 121 17 1697
rect 441 121 475 1697
rect 899 121 933 1697
rect -871 37 -503 71
rect -413 37 -45 71
rect 45 37 413 71
rect 503 37 871 71
rect -933 -1635 -899 -59
rect -475 -1635 -441 -59
rect -17 -1635 17 -59
rect 441 -1635 475 -59
rect 899 -1635 933 -59
rect -871 -1719 -503 -1685
rect -413 -1719 -45 -1685
rect 45 -1719 413 -1685
rect 503 -1719 871 -1685
<< metal1 >>
rect -939 1697 -893 1709
rect -939 121 -933 1697
rect -899 121 -893 1697
rect -939 109 -893 121
rect -481 1697 -435 1709
rect -481 121 -475 1697
rect -441 121 -435 1697
rect -481 109 -435 121
rect -23 1697 23 1709
rect -23 121 -17 1697
rect 17 121 23 1697
rect -23 109 23 121
rect 435 1697 481 1709
rect 435 121 441 1697
rect 475 121 481 1697
rect 435 109 481 121
rect 893 1697 939 1709
rect 893 121 899 1697
rect 933 121 939 1697
rect 893 109 939 121
rect -883 71 -491 77
rect -883 37 -871 71
rect -503 37 -491 71
rect -883 31 -491 37
rect -425 71 -33 77
rect -425 37 -413 71
rect -45 37 -33 71
rect -425 31 -33 37
rect 33 71 425 77
rect 33 37 45 71
rect 413 37 425 71
rect 33 31 425 37
rect 491 71 883 77
rect 491 37 503 71
rect 871 37 883 71
rect 491 31 883 37
rect -939 -59 -893 -47
rect -939 -1635 -933 -59
rect -899 -1635 -893 -59
rect -939 -1647 -893 -1635
rect -481 -59 -435 -47
rect -481 -1635 -475 -59
rect -441 -1635 -435 -59
rect -481 -1647 -435 -1635
rect -23 -59 23 -47
rect -23 -1635 -17 -59
rect 17 -1635 23 -59
rect -23 -1647 23 -1635
rect 435 -59 481 -47
rect 435 -1635 441 -59
rect 475 -1635 481 -59
rect 435 -1647 481 -1635
rect 893 -59 939 -47
rect 893 -1635 899 -59
rect 933 -1635 939 -59
rect 893 -1647 939 -1635
rect -883 -1685 -491 -1679
rect -883 -1719 -871 -1685
rect -503 -1719 -491 -1685
rect -883 -1725 -491 -1719
rect -425 -1685 -33 -1679
rect -425 -1719 -413 -1685
rect -45 -1719 -33 -1685
rect -425 -1725 -33 -1719
rect 33 -1685 425 -1679
rect 33 -1719 45 -1685
rect 413 -1719 425 -1685
rect 33 -1725 425 -1719
rect 491 -1685 883 -1679
rect 491 -1719 503 -1685
rect 871 -1719 883 -1685
rect 491 -1725 883 -1719
<< properties >>
string FIXED_BBOX -1030 -1804 1030 1804
string gencell sky130_fd_pr__nfet_01v8_lvt
string library sky130
string parameters w 8 l 2 m 2 nf 4 diffcov 100 polycov 100 guard 1 glc 0 grc 0 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 0 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
