magic
tech sky130A
magscale 1 2
timestamp 1665771957
<< pwell >>
rect -3223 -11198 3223 11198
<< psubdiff >>
rect -3187 11128 -3091 11162
rect 3091 11128 3187 11162
rect -3187 11066 -3153 11128
rect 3153 11066 3187 11128
rect -3187 -11128 -3153 -11066
rect 3153 -11128 3187 -11066
rect -3187 -11162 -3091 -11128
rect 3091 -11162 3187 -11128
<< psubdiffcont >>
rect -3091 11128 3091 11162
rect -3187 -11066 -3153 11066
rect 3153 -11066 3187 11066
rect -3091 -11162 3091 -11128
<< xpolycontact >>
rect -3057 10600 -1911 11032
rect -3057 -11032 -1911 -10600
rect -1815 10600 -669 11032
rect -1815 -11032 -669 -10600
rect -573 10600 573 11032
rect -573 -11032 573 -10600
rect 669 10600 1815 11032
rect 669 -11032 1815 -10600
rect 1911 10600 3057 11032
rect 1911 -11032 3057 -10600
<< xpolyres >>
rect -3057 -10600 -1911 10600
rect -1815 -10600 -669 10600
rect -573 -10600 573 10600
rect 669 -10600 1815 10600
rect 1911 -10600 3057 10600
<< locali >>
rect -3187 11128 -3091 11162
rect 3091 11128 3187 11162
rect -3187 11066 -3153 11128
rect 3153 11066 3187 11128
rect -3187 -11128 -3153 -11066
rect 3153 -11128 3187 -11066
rect -3187 -11162 -3091 -11128
rect 3091 -11162 3187 -11128
<< viali >>
rect -3041 10617 -1927 11014
rect -1799 10617 -685 11014
rect -557 10617 557 11014
rect 685 10617 1799 11014
rect 1927 10617 3041 11014
rect -3041 -11014 -1927 -10617
rect -1799 -11014 -685 -10617
rect -557 -11014 557 -10617
rect 685 -11014 1799 -10617
rect 1927 -11014 3041 -10617
<< metal1 >>
rect -3053 11014 -1915 11020
rect -3053 10617 -3041 11014
rect -1927 10617 -1915 11014
rect -3053 10611 -1915 10617
rect -1811 11014 -673 11020
rect -1811 10617 -1799 11014
rect -685 10617 -673 11014
rect -1811 10611 -673 10617
rect -569 11014 569 11020
rect -569 10617 -557 11014
rect 557 10617 569 11014
rect -569 10611 569 10617
rect 673 11014 1811 11020
rect 673 10617 685 11014
rect 1799 10617 1811 11014
rect 673 10611 1811 10617
rect 1915 11014 3053 11020
rect 1915 10617 1927 11014
rect 3041 10617 3053 11014
rect 1915 10611 3053 10617
rect -3053 -10617 -1915 -10611
rect -3053 -11014 -3041 -10617
rect -1927 -11014 -1915 -10617
rect -3053 -11020 -1915 -11014
rect -1811 -10617 -673 -10611
rect -1811 -11014 -1799 -10617
rect -685 -11014 -673 -10617
rect -1811 -11020 -673 -11014
rect -569 -10617 569 -10611
rect -569 -11014 -557 -10617
rect 557 -11014 569 -10617
rect -569 -11020 569 -11014
rect 673 -10617 1811 -10611
rect 673 -11014 685 -10617
rect 1799 -11014 1811 -10617
rect 673 -11020 1811 -11014
rect 1915 -10617 3053 -10611
rect 1915 -11014 1927 -10617
rect 3041 -11014 3053 -10617
rect 1915 -11020 3053 -11014
<< res5p73 >>
rect -3059 -10602 -1909 10602
rect -1817 -10602 -667 10602
rect -575 -10602 575 10602
rect 667 -10602 1817 10602
rect 1909 -10602 3059 10602
<< properties >>
string FIXED_BBOX -3170 -11145 3170 11145
string gencell sky130_fd_pr__res_xhigh_po_5p73
string library sky130
string parameters w 5.730 l 106 m 1 nx 5 wmin 5.730 lmin 0.50 rho 2000 val 37.063k dummy 0 dw 0.0 term 188.2 sterm 0.0 caplen 0 wmax 5.730 guard 1 glc 1 grc 1 gtc 1 gbc 1 compatible {sky130_fd_pr__res_xhigh_po_0p35  sky130_fd_pr__res_xhigh_po_0p69 sky130_fd_pr__res_xhigh_po_1p41  sky130_fd_pr__res_xhigh_po_2p85 sky130_fd_pr__res_xhigh_po_5p73} snake 0 full_metal 1 n_guard 0 hv_guard 0 vias 1 viagb 0 viagt 0 viagl 0 viagr 0
<< end >>
