magic
tech sky130A
magscale 1 2
timestamp 1662517639
<< pwell >>
rect 14375 550 14421 750
rect 14565 550 14611 750
rect 14665 550 14711 750
rect 14760 550 14806 750
rect 14855 550 14901 750
rect 14950 550 14996 750
rect 15050 550 15096 750
rect 15145 550 15191 750
rect 15240 550 15286 750
rect 15335 550 15381 750
rect 15430 550 15476 750
rect 15525 550 15571 750
rect 15625 550 15671 750
rect 16385 550 16430 750
rect 16485 550 16530 750
rect 16580 550 16625 750
rect 16675 550 16720 750
rect 16770 550 16815 750
rect 16870 550 16915 750
rect 16965 550 17010 750
rect 17060 550 17105 750
rect 17155 550 17200 750
rect 17250 550 17295 750
rect 17350 550 17395 750
rect 17445 550 17490 750
rect 17540 550 17585 750
rect 17635 550 17680 750
rect 17735 550 17780 750
rect 17830 550 17875 750
rect 17925 550 17970 750
rect 18020 550 18065 750
rect 18115 550 18160 750
rect 18210 550 18255 750
rect 18310 550 18355 750
rect 18405 550 18450 750
rect 18500 550 18545 750
rect 18690 550 18735 750
rect 18790 550 18835 750
rect 18885 550 18930 750
rect 18980 550 19025 750
rect 19075 550 19120 750
rect 19170 550 19215 750
rect 19270 550 19315 750
rect 19365 550 19410 750
rect 19460 550 19505 750
rect 19555 550 19600 750
rect 19650 550 19695 750
rect 19750 550 19795 750
rect 19845 550 19890 750
rect 19940 550 19985 750
rect 20035 550 20080 750
rect 20135 550 20180 750
rect 20230 550 20275 750
rect 20325 550 20370 750
rect 20420 550 20465 750
rect 20515 550 20560 750
rect 20610 550 20655 750
rect 20710 550 20755 750
rect 20805 550 20850 750
rect 20900 550 20945 750
rect 20995 550 21040 750
rect 21090 550 21135 750
rect 21190 550 21235 750
rect 21285 550 21330 750
rect 21380 550 21425 750
rect 21475 550 21520 750
rect 21570 550 21615 750
rect 21670 550 21715 750
rect 21765 550 21810 750
<< ndiff >>
rect 14375 550 14421 750
<< locali >>
rect 12675 1830 13610 1870
rect 10060 880 10095 1110
rect 12665 1070 13615 1075
rect 11900 925 11935 1070
rect 12055 925 12090 1070
rect 11900 885 12090 925
rect 12665 1035 13630 1070
rect 12665 930 12705 1035
rect 13595 930 13630 1035
rect 12665 890 13630 930
rect 15745 920 15780 1075
rect 15895 920 15930 1070
rect 15745 890 15930 920
rect 17960 890 17995 1140
rect 12665 885 12705 890
rect 15745 885 15925 890
rect 9755 230 9795 420
rect 11905 235 11945 425
rect 12050 230 12090 420
rect 12690 415 13625 420
rect 12665 405 13625 415
rect 12665 380 13635 405
rect 12665 265 12705 380
rect 13600 265 13635 380
rect 12665 225 13635 265
rect 15735 230 15770 410
rect 15910 230 15945 410
rect 21885 225 21920 415
rect 11905 -250 12090 -245
rect 10055 -430 10095 -250
rect 11905 -285 12095 -250
rect 11905 -430 11945 -285
rect 12055 -430 12095 -285
rect 12660 -260 13625 -250
rect 15740 -255 15775 -245
rect 15895 -255 15930 -245
rect 12660 -290 13630 -260
rect 12660 -400 12700 -290
rect 13595 -400 13630 -290
rect 12660 -430 13630 -400
rect 15740 -290 15930 -255
rect 15740 -425 15775 -290
rect 15895 -425 15930 -290
rect 12680 -440 13630 -430
rect 17965 -435 18005 -250
rect 12675 -1220 13610 -1180
<< metal1 >>
rect 17435 2280 17870 2310
rect 12140 1720 12590 1735
rect 12140 1185 12170 1720
rect 12575 1185 12590 1720
rect 17435 1190 17455 2280
rect 17840 1190 17870 2280
rect 12140 1165 12590 1185
rect 17435 1165 17870 1190
rect 13515 850 13590 860
rect 9900 780 11975 830
rect 12190 780 12740 830
rect 13515 795 13525 850
rect 13580 835 13590 850
rect 13580 795 15675 835
rect 13515 785 15675 795
rect 9860 625 9910 750
rect 9945 740 10020 750
rect 9945 685 9955 740
rect 10010 685 10020 740
rect 9945 675 10020 685
rect 9850 615 9925 625
rect 9850 560 9860 615
rect 9915 560 9925 615
rect 9850 550 9925 560
rect 9960 550 10010 675
rect 10050 625 10100 750
rect 10140 740 10215 750
rect 10140 685 10150 740
rect 10205 685 10215 740
rect 10140 675 10215 685
rect 10040 615 10115 625
rect 10040 560 10050 615
rect 10105 560 10115 615
rect 10040 550 10115 560
rect 10150 550 10200 675
rect 10250 625 10300 750
rect 10330 740 10405 750
rect 10330 685 10340 740
rect 10395 685 10405 740
rect 10330 675 10405 685
rect 10230 615 10305 625
rect 10230 560 10240 615
rect 10295 560 10305 615
rect 10230 550 10305 560
rect 10340 550 10390 675
rect 10440 625 10490 750
rect 10520 740 10595 750
rect 10520 685 10530 740
rect 10585 685 10595 740
rect 10520 675 10595 685
rect 10420 615 10495 625
rect 10420 560 10430 615
rect 10485 560 10495 615
rect 10420 550 10495 560
rect 10530 550 10580 675
rect 10630 625 10680 750
rect 10710 740 10785 750
rect 10710 685 10720 740
rect 10775 685 10785 740
rect 10710 675 10785 685
rect 10620 615 10695 625
rect 10620 560 10630 615
rect 10685 560 10695 615
rect 10620 550 10695 560
rect 10730 550 10780 675
rect 10820 625 10870 750
rect 10900 740 10975 750
rect 10900 685 10910 740
rect 10965 685 10975 740
rect 10900 675 10975 685
rect 10810 615 10885 625
rect 10810 560 10820 615
rect 10875 560 10885 615
rect 10810 550 10885 560
rect 10920 550 10970 675
rect 11010 625 11060 750
rect 11095 740 11170 750
rect 11095 685 11105 740
rect 11160 685 11170 740
rect 11095 675 11170 685
rect 11005 615 11080 625
rect 11005 560 11015 615
rect 11070 560 11080 615
rect 11005 550 11080 560
rect 11110 550 11160 675
rect 11210 625 11260 750
rect 11290 740 11365 750
rect 11290 685 11300 740
rect 11355 685 11365 740
rect 11290 675 11365 685
rect 11195 615 11270 625
rect 11195 560 11205 615
rect 11260 560 11270 615
rect 11195 550 11270 560
rect 11300 550 11350 675
rect 11400 625 11450 750
rect 11480 740 11555 750
rect 11480 685 11490 740
rect 11545 685 11555 740
rect 11480 675 11555 685
rect 11385 615 11460 625
rect 11385 560 11395 615
rect 11450 560 11460 615
rect 11385 550 11460 560
rect 11490 550 11540 675
rect 11590 625 11640 750
rect 11675 740 11750 750
rect 11675 685 11685 740
rect 11740 685 11750 740
rect 11675 675 11750 685
rect 11580 615 11655 625
rect 11580 560 11590 615
rect 11645 560 11655 615
rect 11580 550 11655 560
rect 11690 550 11740 675
rect 11780 625 11830 750
rect 11770 615 11845 625
rect 11770 560 11780 615
rect 11835 560 11845 615
rect 11770 550 11845 560
rect 11925 520 11975 780
rect 12165 625 12215 750
rect 12245 740 12320 750
rect 12245 685 12255 740
rect 12310 685 12320 740
rect 12245 675 12320 685
rect 12150 615 12225 625
rect 12150 560 12160 615
rect 12215 560 12225 615
rect 12150 550 12225 560
rect 12255 550 12306 675
rect 12350 625 12401 750
rect 12435 740 12510 750
rect 12435 685 12445 740
rect 12500 685 12510 740
rect 12435 675 12510 685
rect 12340 615 12415 625
rect 12340 560 12350 615
rect 12405 560 12415 615
rect 12340 550 12415 560
rect 12450 550 12501 675
rect 12545 625 12596 750
rect 12535 615 12610 625
rect 12535 560 12545 615
rect 12600 560 12610 615
rect 12535 550 12610 560
rect 12685 520 12740 780
rect 13535 520 13585 785
rect 15855 780 21775 830
rect 13785 740 13860 750
rect 13785 685 13795 740
rect 13850 685 13860 740
rect 13785 675 13860 685
rect 13705 625 13750 670
rect 13690 615 13765 625
rect 13690 560 13700 615
rect 13755 560 13765 615
rect 13690 550 13765 560
rect 13800 550 13846 675
rect 13895 625 13941 750
rect 13975 740 14050 750
rect 13975 685 13985 740
rect 14040 685 14050 740
rect 13975 675 14050 685
rect 13880 615 13955 625
rect 13880 560 13890 615
rect 13945 560 13955 615
rect 13880 550 13955 560
rect 13990 550 14036 675
rect 14085 625 14131 750
rect 14170 740 14245 750
rect 14170 685 14180 740
rect 14235 685 14245 740
rect 14170 675 14245 685
rect 14075 615 14150 625
rect 14075 560 14085 615
rect 14140 560 14150 615
rect 14075 550 14150 560
rect 14185 550 14231 675
rect 14280 625 14326 750
rect 14360 740 14435 750
rect 14360 685 14370 740
rect 14425 685 14435 740
rect 14360 675 14435 685
rect 14265 615 14340 625
rect 14265 560 14275 615
rect 14330 560 14340 615
rect 14265 550 14340 560
rect 14375 550 14421 675
rect 14470 625 14516 750
rect 14550 740 14625 750
rect 14550 685 14560 740
rect 14615 685 14625 740
rect 14550 675 14625 685
rect 14460 615 14535 625
rect 14460 560 14470 615
rect 14525 560 14535 615
rect 14460 550 14535 560
rect 14565 550 14611 675
rect 14665 625 14711 750
rect 14745 740 14820 750
rect 14745 685 14755 740
rect 14810 685 14820 740
rect 14745 675 14820 685
rect 14645 615 14720 625
rect 14645 560 14655 615
rect 14710 560 14720 615
rect 14645 550 14720 560
rect 14760 550 14806 675
rect 14855 625 14901 750
rect 14935 740 15010 750
rect 14935 685 14945 740
rect 15000 685 15010 740
rect 14935 675 15010 685
rect 14840 615 14915 625
rect 14840 560 14850 615
rect 14905 560 14915 615
rect 14840 550 14915 560
rect 14950 550 14996 675
rect 15050 625 15096 750
rect 15130 740 15205 750
rect 15130 685 15140 740
rect 15195 685 15205 740
rect 15130 675 15205 685
rect 15030 615 15105 625
rect 15030 560 15040 615
rect 15095 560 15105 615
rect 15030 550 15105 560
rect 15145 550 15191 675
rect 15240 625 15286 750
rect 15320 740 15395 750
rect 15320 685 15330 740
rect 15385 685 15395 740
rect 15320 675 15395 685
rect 15225 615 15300 625
rect 15225 560 15235 615
rect 15290 560 15300 615
rect 15225 550 15300 560
rect 15335 550 15381 675
rect 15430 625 15476 750
rect 15510 740 15585 750
rect 15510 685 15520 740
rect 15575 685 15585 740
rect 15510 675 15585 685
rect 15415 615 15490 625
rect 15415 560 15425 615
rect 15480 560 15490 615
rect 15415 550 15490 560
rect 15525 550 15571 675
rect 15625 625 15671 750
rect 15610 615 15685 625
rect 15610 560 15620 615
rect 15675 560 15685 615
rect 15610 550 15685 560
rect 9990 470 11975 520
rect 12295 470 13415 520
rect 13535 470 15625 520
rect 15855 515 15905 780
rect 16005 625 16050 750
rect 16085 740 16160 750
rect 16085 685 16095 740
rect 16150 685 16160 740
rect 16085 675 16160 685
rect 15985 615 16060 625
rect 15985 560 15995 615
rect 16050 560 16060 615
rect 15985 550 16060 560
rect 16100 550 16145 675
rect 16195 625 16240 750
rect 16275 740 16350 750
rect 16275 685 16285 740
rect 16340 685 16350 740
rect 16275 675 16350 685
rect 16175 615 16250 625
rect 16175 560 16185 615
rect 16240 560 16250 615
rect 16175 550 16250 560
rect 16290 550 16335 675
rect 16385 625 16430 750
rect 16470 740 16545 750
rect 16470 685 16480 740
rect 16535 685 16545 740
rect 16470 675 16545 685
rect 16370 615 16445 625
rect 16370 560 16380 615
rect 16435 560 16445 615
rect 16370 550 16445 560
rect 16485 550 16530 675
rect 16580 625 16625 750
rect 16660 740 16735 750
rect 16660 685 16670 740
rect 16725 685 16735 740
rect 16660 675 16735 685
rect 16565 615 16640 625
rect 16565 560 16575 615
rect 16630 560 16640 615
rect 16565 550 16640 560
rect 16675 550 16720 675
rect 16770 625 16815 750
rect 16855 740 16930 750
rect 16855 685 16865 740
rect 16920 685 16930 740
rect 16855 675 16930 685
rect 16755 615 16830 625
rect 16755 560 16765 615
rect 16820 560 16830 615
rect 16755 550 16830 560
rect 16870 550 16915 675
rect 16965 625 17010 750
rect 17040 740 17115 750
rect 17040 685 17050 740
rect 17105 685 17115 740
rect 17040 675 17115 685
rect 16950 615 17025 625
rect 16950 560 16960 615
rect 17015 560 17025 615
rect 16950 550 17025 560
rect 17060 550 17105 675
rect 17155 625 17200 750
rect 17240 740 17315 750
rect 17240 685 17250 740
rect 17305 685 17315 740
rect 17240 675 17315 685
rect 17140 615 17215 625
rect 17140 560 17150 615
rect 17205 560 17215 615
rect 17140 550 17215 560
rect 17250 550 17295 675
rect 17350 625 17395 750
rect 17425 740 17500 750
rect 17425 685 17435 740
rect 17490 685 17500 740
rect 17425 675 17500 685
rect 17335 615 17410 625
rect 17335 560 17345 615
rect 17400 560 17410 615
rect 17335 550 17410 560
rect 17445 550 17490 675
rect 17540 625 17585 750
rect 17620 740 17695 750
rect 17620 685 17630 740
rect 17685 685 17695 740
rect 17620 675 17695 685
rect 17525 615 17600 625
rect 17525 560 17535 615
rect 17590 560 17600 615
rect 17525 550 17600 560
rect 17635 550 17680 675
rect 17735 625 17780 750
rect 17815 740 17890 750
rect 17815 685 17825 740
rect 17880 685 17890 740
rect 17815 675 17890 685
rect 17715 615 17790 625
rect 17715 560 17725 615
rect 17780 560 17790 615
rect 17715 550 17790 560
rect 17830 550 17875 675
rect 17925 625 17970 750
rect 18000 740 18075 750
rect 18000 685 18010 740
rect 18065 685 18075 740
rect 18000 675 18075 685
rect 17910 615 17985 625
rect 17910 560 17920 615
rect 17975 560 17985 615
rect 17910 550 17985 560
rect 18020 550 18065 675
rect 18115 625 18160 750
rect 18195 740 18270 750
rect 18195 685 18205 740
rect 18260 685 18270 740
rect 18195 675 18270 685
rect 18100 615 18175 625
rect 18100 560 18110 615
rect 18165 560 18175 615
rect 18100 550 18175 560
rect 18210 550 18255 675
rect 18310 625 18355 750
rect 18385 740 18460 750
rect 18385 685 18395 740
rect 18450 685 18460 740
rect 18385 675 18460 685
rect 18295 615 18370 625
rect 18295 560 18305 615
rect 18360 560 18370 615
rect 18295 550 18370 560
rect 18405 550 18450 675
rect 18500 625 18545 750
rect 18580 740 18655 750
rect 18580 685 18590 740
rect 18645 685 18655 740
rect 18580 675 18655 685
rect 18485 615 18560 625
rect 18485 560 18495 615
rect 18550 560 18560 615
rect 18485 550 18560 560
rect 18595 550 18640 675
rect 18690 625 18735 750
rect 18770 740 18845 750
rect 18770 685 18780 740
rect 18835 685 18845 740
rect 18770 675 18845 685
rect 18675 615 18750 625
rect 18675 560 18685 615
rect 18740 560 18750 615
rect 18675 550 18750 560
rect 18790 550 18835 675
rect 18885 625 18930 750
rect 18965 740 19040 750
rect 18965 685 18975 740
rect 19030 685 19040 740
rect 18965 675 19040 685
rect 18870 615 18945 625
rect 18870 560 18880 615
rect 18935 560 18945 615
rect 18870 550 18945 560
rect 18980 550 19025 675
rect 19075 625 19120 750
rect 19155 740 19230 750
rect 19155 685 19165 740
rect 19220 685 19230 740
rect 19155 675 19230 685
rect 19060 615 19135 625
rect 19060 560 19070 615
rect 19125 560 19135 615
rect 19060 550 19135 560
rect 19170 550 19215 675
rect 19270 625 19315 750
rect 19350 740 19425 750
rect 19350 685 19360 740
rect 19415 685 19425 740
rect 19350 675 19425 685
rect 19255 615 19330 625
rect 19255 560 19265 615
rect 19320 560 19330 615
rect 19255 550 19330 560
rect 19365 550 19410 675
rect 19460 625 19505 750
rect 19540 740 19615 750
rect 19540 685 19550 740
rect 19605 685 19615 740
rect 19540 675 19615 685
rect 19445 615 19520 625
rect 19445 560 19455 615
rect 19510 560 19520 615
rect 19445 550 19520 560
rect 19555 550 19600 675
rect 19650 625 19695 750
rect 19735 740 19810 750
rect 19735 685 19745 740
rect 19800 685 19810 740
rect 19735 675 19810 685
rect 19635 615 19710 625
rect 19635 560 19645 615
rect 19700 560 19710 615
rect 19635 550 19710 560
rect 19750 550 19795 675
rect 19845 625 19890 750
rect 19925 740 20000 750
rect 19925 685 19935 740
rect 19990 685 20000 740
rect 19925 675 20000 685
rect 19830 615 19905 625
rect 19830 560 19840 615
rect 19895 560 19905 615
rect 19830 550 19905 560
rect 19940 550 19985 675
rect 20035 625 20080 750
rect 20115 740 20190 750
rect 20115 685 20125 740
rect 20180 685 20190 740
rect 20115 675 20190 685
rect 20020 615 20095 625
rect 20020 560 20030 615
rect 20085 560 20095 615
rect 20020 550 20095 560
rect 20135 550 20180 675
rect 20230 625 20275 750
rect 20310 740 20385 750
rect 20310 685 20320 740
rect 20375 685 20385 740
rect 20310 675 20385 685
rect 20215 615 20290 625
rect 20215 560 20225 615
rect 20280 560 20290 615
rect 20215 550 20290 560
rect 20325 550 20370 675
rect 20420 625 20465 750
rect 20500 740 20575 750
rect 20500 685 20510 740
rect 20565 685 20575 740
rect 20500 675 20575 685
rect 20405 615 20480 625
rect 20405 560 20415 615
rect 20470 560 20480 615
rect 20405 550 20480 560
rect 20515 550 20560 675
rect 20610 625 20655 750
rect 20695 740 20770 750
rect 20695 685 20705 740
rect 20760 685 20770 740
rect 20695 675 20770 685
rect 20600 615 20675 625
rect 20600 560 20610 615
rect 20665 560 20675 615
rect 20600 550 20675 560
rect 20710 550 20755 675
rect 20805 625 20850 750
rect 20885 740 20960 750
rect 20885 685 20895 740
rect 20950 685 20960 740
rect 20885 675 20960 685
rect 20790 615 20865 625
rect 20790 560 20800 615
rect 20855 560 20865 615
rect 20790 550 20865 560
rect 20900 550 20945 675
rect 20995 625 21040 750
rect 21075 740 21150 750
rect 21075 685 21085 740
rect 21140 685 21150 740
rect 21075 675 21150 685
rect 20980 615 21055 625
rect 20980 560 20990 615
rect 21045 560 21055 615
rect 20980 550 21055 560
rect 21090 550 21135 675
rect 21190 625 21235 750
rect 21270 740 21345 750
rect 21270 685 21280 740
rect 21335 685 21345 740
rect 21270 675 21345 685
rect 21175 615 21250 625
rect 21175 560 21185 615
rect 21240 560 21250 615
rect 21175 550 21250 560
rect 21285 550 21330 675
rect 21380 625 21425 750
rect 21460 740 21535 750
rect 21460 685 21470 740
rect 21525 685 21535 740
rect 21460 675 21535 685
rect 21365 615 21440 625
rect 21365 560 21375 615
rect 21430 560 21440 615
rect 21365 550 21440 560
rect 21475 550 21520 675
rect 21570 625 21615 750
rect 21650 740 21725 750
rect 21650 685 21660 740
rect 21715 685 21725 740
rect 21650 675 21725 685
rect 21555 615 21630 625
rect 21555 560 21565 615
rect 21620 560 21630 615
rect 21555 550 21630 560
rect 21670 550 21715 675
rect 21765 625 21810 750
rect 21750 615 21825 625
rect 21750 560 21760 615
rect 21815 560 21825 615
rect 21750 550 21825 560
rect 11925 170 11975 470
rect 9990 120 11975 170
rect 12290 125 12955 175
rect 12295 120 12955 125
rect 9850 80 9925 90
rect 9850 25 9860 80
rect 9915 25 9925 80
rect 9850 15 9925 25
rect 9860 -110 9910 15
rect 9960 -35 10010 90
rect 10040 80 10115 90
rect 10040 25 10050 80
rect 10105 25 10115 80
rect 10040 15 10115 25
rect 9945 -45 10020 -35
rect 9945 -100 9955 -45
rect 10010 -100 10020 -45
rect 9945 -110 10020 -100
rect 10050 -110 10102 15
rect 10150 -35 10200 90
rect 10230 80 10305 90
rect 10230 25 10240 80
rect 10295 25 10305 80
rect 10230 15 10305 25
rect 10140 -45 10215 -35
rect 10140 -100 10150 -45
rect 10205 -100 10215 -45
rect 10140 -110 10215 -100
rect 10248 -110 10300 15
rect 10340 -35 10390 90
rect 10420 80 10495 90
rect 10420 25 10430 80
rect 10485 25 10495 80
rect 10420 15 10495 25
rect 10330 -45 10405 -35
rect 10330 -100 10340 -45
rect 10395 -100 10405 -45
rect 10330 -110 10405 -100
rect 10440 -110 10490 15
rect 10530 -35 10582 90
rect 10620 80 10695 90
rect 10620 25 10630 80
rect 10685 25 10695 80
rect 10620 15 10695 25
rect 10520 -45 10595 -35
rect 10520 -100 10530 -45
rect 10585 -100 10595 -45
rect 10520 -110 10595 -100
rect 10630 -110 10680 15
rect 10728 -35 10780 90
rect 10810 80 10885 90
rect 10810 25 10820 80
rect 10875 25 10885 80
rect 10810 15 10885 25
rect 10710 -45 10785 -35
rect 10710 -100 10720 -45
rect 10775 -100 10785 -45
rect 10710 -110 10785 -100
rect 10820 -110 10870 15
rect 10920 -35 10970 90
rect 11005 80 11080 90
rect 11005 25 11015 80
rect 11070 25 11080 80
rect 11005 15 11080 25
rect 10900 -45 10975 -35
rect 10900 -100 10910 -45
rect 10965 -100 10975 -45
rect 10900 -110 10975 -100
rect 11010 -110 11062 15
rect 11110 -35 11160 90
rect 11195 80 11270 90
rect 11195 25 11205 80
rect 11260 25 11270 80
rect 11195 15 11270 25
rect 11095 -45 11170 -35
rect 11095 -100 11105 -45
rect 11160 -100 11170 -45
rect 11095 -110 11170 -100
rect 11208 -110 11260 15
rect 11300 -35 11350 90
rect 11385 80 11460 90
rect 11385 25 11395 80
rect 11450 25 11460 80
rect 11385 15 11460 25
rect 11290 -45 11365 -35
rect 11290 -100 11300 -45
rect 11355 -100 11365 -45
rect 11290 -110 11365 -100
rect 11400 -110 11450 15
rect 11490 -35 11542 90
rect 11580 80 11655 90
rect 11580 25 11590 80
rect 11645 25 11655 80
rect 11580 15 11655 25
rect 11480 -45 11555 -35
rect 11480 -100 11490 -45
rect 11545 -100 11555 -45
rect 11480 -110 11555 -100
rect 11590 -110 11640 15
rect 11688 -35 11740 90
rect 11770 80 11845 90
rect 11770 25 11780 80
rect 11835 25 11845 80
rect 11770 15 11845 25
rect 11675 -45 11750 -35
rect 11675 -100 11685 -45
rect 11740 -100 11750 -45
rect 11675 -110 11750 -100
rect 11780 -110 11830 15
rect 11925 -140 11975 120
rect 12150 80 12225 90
rect 12150 25 12160 80
rect 12215 25 12225 80
rect 12150 15 12225 25
rect 12164 -110 12215 15
rect 12255 -35 12306 90
rect 12340 80 12415 90
rect 12340 25 12350 80
rect 12405 25 12415 80
rect 12340 15 12415 25
rect 12245 -45 12320 -35
rect 12245 -100 12255 -45
rect 12310 -100 12320 -45
rect 12245 -110 12320 -100
rect 12350 -110 12402 15
rect 12450 -35 12501 90
rect 12535 80 12610 90
rect 12535 25 12545 80
rect 12600 25 12610 80
rect 12535 15 12610 25
rect 12435 -45 12510 -35
rect 12435 -100 12445 -45
rect 12500 -100 12510 -45
rect 12435 -110 12510 -100
rect 12545 -110 12596 15
rect 12685 -140 12740 120
rect 9900 -190 11975 -140
rect 12190 -190 12740 -140
rect 11925 -1260 11975 -190
rect 12200 -195 12740 -190
rect 12140 -540 12570 -525
rect 12140 -1075 12160 -540
rect 12550 -1075 12570 -540
rect 12140 -1090 12570 -1075
rect 12900 -1255 12955 120
rect 13365 -1260 13415 470
rect 15855 465 21775 515
rect 15855 175 15905 465
rect 13535 120 15625 170
rect 15855 125 21775 175
rect 13535 -145 13585 120
rect 13690 80 13765 90
rect 13690 25 13700 80
rect 13755 25 13765 80
rect 13690 15 13765 25
rect 13704 -30 13750 15
rect 13704 -98 13710 -30
rect 13744 -98 13750 -30
rect 13800 -35 13846 90
rect 13880 80 13955 90
rect 13880 25 13890 80
rect 13945 25 13955 80
rect 13880 15 13955 25
rect 13704 -110 13750 -98
rect 13785 -45 13860 -35
rect 13785 -100 13795 -45
rect 13850 -100 13860 -45
rect 13785 -110 13860 -100
rect 13895 -110 13942 15
rect 13990 -35 14038 90
rect 14075 80 14150 90
rect 14075 25 14085 80
rect 14140 25 14150 80
rect 14075 15 14150 25
rect 13975 -45 14050 -35
rect 13975 -100 13985 -45
rect 14040 -100 14050 -45
rect 13975 -110 14050 -100
rect 14085 -110 14134 15
rect 14184 -35 14231 90
rect 14265 80 14340 90
rect 14265 25 14275 80
rect 14330 25 14340 80
rect 14265 15 14340 25
rect 14170 -45 14245 -35
rect 14170 -100 14180 -45
rect 14235 -100 14245 -45
rect 14170 -110 14245 -100
rect 14280 -110 14326 15
rect 14375 -35 14422 90
rect 14460 80 14535 90
rect 14460 25 14470 80
rect 14525 25 14535 80
rect 14460 15 14535 25
rect 14360 -45 14435 -35
rect 14360 -100 14370 -45
rect 14425 -100 14435 -45
rect 14360 -110 14435 -100
rect 14470 -110 14518 15
rect 14565 -35 14614 90
rect 14645 80 14720 90
rect 14645 25 14655 80
rect 14710 25 14720 80
rect 14645 15 14720 25
rect 14550 -45 14625 -35
rect 14550 -100 14560 -45
rect 14615 -100 14625 -45
rect 14550 -110 14625 -100
rect 14664 -110 14711 15
rect 14760 -35 14806 90
rect 14840 80 14915 90
rect 14840 25 14850 80
rect 14905 25 14915 80
rect 14840 15 14915 25
rect 14745 -45 14820 -35
rect 14745 -100 14755 -45
rect 14810 -100 14820 -45
rect 14745 -110 14820 -100
rect 14855 -110 14902 15
rect 14950 -35 14998 90
rect 15030 80 15105 90
rect 15030 25 15040 80
rect 15095 25 15105 80
rect 15030 15 15105 25
rect 14935 -45 15010 -35
rect 14935 -100 14945 -45
rect 15000 -100 15010 -45
rect 14935 -110 15010 -100
rect 15048 -110 15096 15
rect 15144 -35 15191 90
rect 15225 80 15300 90
rect 15225 25 15235 80
rect 15290 25 15300 80
rect 15225 15 15300 25
rect 15130 -45 15205 -35
rect 15130 -100 15140 -45
rect 15195 -100 15205 -45
rect 15130 -110 15205 -100
rect 15240 -110 15286 15
rect 15335 -35 15382 90
rect 15415 80 15490 90
rect 15415 25 15425 80
rect 15480 25 15490 80
rect 15415 15 15490 25
rect 15320 -45 15395 -35
rect 15320 -100 15330 -45
rect 15385 -100 15395 -45
rect 15320 -110 15395 -100
rect 15430 -110 15478 15
rect 15525 -35 15574 90
rect 15610 80 15685 90
rect 15610 25 15620 80
rect 15675 25 15685 80
rect 15610 15 15685 25
rect 15510 -45 15585 -35
rect 15510 -100 15520 -45
rect 15575 -100 15585 -45
rect 15510 -110 15585 -100
rect 15624 -110 15671 15
rect 15855 -140 15905 125
rect 16046 122 16104 125
rect 16238 122 16296 125
rect 16430 122 16488 125
rect 16622 122 16680 125
rect 16814 122 16872 125
rect 17006 122 17064 125
rect 17198 122 17256 125
rect 17390 122 17448 125
rect 17582 122 17640 125
rect 17774 122 17832 125
rect 17966 122 18024 125
rect 18158 122 18216 125
rect 18350 122 18408 125
rect 18542 122 18600 125
rect 18734 122 18792 125
rect 18926 122 18984 125
rect 19118 122 19176 125
rect 19310 122 19368 125
rect 19502 122 19560 125
rect 19694 122 19752 125
rect 19886 122 19944 125
rect 20078 122 20136 125
rect 20270 122 20328 125
rect 20462 122 20520 125
rect 20654 122 20712 125
rect 20846 122 20904 125
rect 21038 122 21096 125
rect 21230 122 21288 125
rect 21422 122 21480 125
rect 21614 122 21672 125
rect 15985 80 16060 90
rect 15985 25 15995 80
rect 16050 25 16060 80
rect 15985 15 16060 25
rect 16004 -110 16050 15
rect 16100 -35 16146 90
rect 16175 80 16250 90
rect 16175 25 16185 80
rect 16240 25 16250 80
rect 16175 15 16250 25
rect 16085 -45 16160 -35
rect 16085 -100 16095 -45
rect 16150 -100 16160 -45
rect 16085 -110 16160 -100
rect 16195 -110 16242 15
rect 16290 -35 16338 90
rect 16370 80 16445 90
rect 16370 25 16380 80
rect 16435 25 16445 80
rect 16370 15 16445 25
rect 16275 -45 16350 -35
rect 16275 -100 16285 -45
rect 16340 -100 16350 -45
rect 16275 -110 16350 -100
rect 16385 -110 16434 15
rect 16484 -35 16530 90
rect 16565 80 16640 90
rect 16565 25 16575 80
rect 16630 25 16640 80
rect 16565 15 16640 25
rect 16470 -45 16545 -35
rect 16470 -100 16480 -45
rect 16535 -100 16545 -45
rect 16470 -110 16545 -100
rect 16580 -110 16626 15
rect 16675 -35 16722 90
rect 16755 80 16830 90
rect 16755 25 16765 80
rect 16820 25 16830 80
rect 16755 15 16830 25
rect 16660 -45 16735 -35
rect 16660 -100 16670 -45
rect 16725 -100 16735 -45
rect 16660 -110 16735 -100
rect 16770 -110 16818 15
rect 16868 -35 16915 90
rect 16950 80 17025 90
rect 16950 25 16960 80
rect 17015 25 17025 80
rect 16950 15 17025 25
rect 16855 -45 16930 -35
rect 16855 -100 16865 -45
rect 16920 -100 16930 -45
rect 16855 -110 16930 -100
rect 16964 -110 17010 15
rect 17060 -35 17106 90
rect 17140 80 17215 90
rect 17140 25 17150 80
rect 17205 25 17215 80
rect 17140 15 17215 25
rect 17040 -45 17115 -35
rect 17040 -100 17050 -45
rect 17105 -100 17115 -45
rect 17040 -110 17115 -100
rect 17155 -110 17202 15
rect 17250 -35 17298 90
rect 17335 80 17410 90
rect 17335 25 17345 80
rect 17400 25 17410 80
rect 17335 15 17410 25
rect 17240 -45 17315 -35
rect 17240 -100 17250 -45
rect 17305 -100 17315 -45
rect 17240 -110 17315 -100
rect 17348 -110 17395 15
rect 17444 -35 17490 90
rect 17525 80 17600 90
rect 17525 25 17535 80
rect 17590 25 17600 80
rect 17525 15 17600 25
rect 17425 -45 17500 -35
rect 17425 -100 17435 -45
rect 17490 -100 17500 -45
rect 17425 -110 17500 -100
rect 17540 -110 17586 15
rect 17635 -35 17682 90
rect 17715 80 17790 90
rect 17715 25 17725 80
rect 17780 25 17790 80
rect 17715 15 17790 25
rect 17620 -45 17695 -35
rect 17620 -100 17630 -45
rect 17685 -100 17695 -45
rect 17620 -110 17695 -100
rect 17732 -110 17780 15
rect 17828 -35 17875 90
rect 17910 80 17985 90
rect 17910 25 17920 80
rect 17975 25 17985 80
rect 17910 15 17985 25
rect 17815 -45 17890 -35
rect 17815 -100 17825 -45
rect 17880 -100 17890 -45
rect 17815 -110 17890 -100
rect 17924 -110 17970 15
rect 18020 -35 18066 90
rect 18100 80 18175 90
rect 18100 25 18110 80
rect 18165 25 18175 80
rect 18100 15 18175 25
rect 18000 -45 18075 -35
rect 18000 -100 18010 -45
rect 18065 -100 18075 -45
rect 18000 -110 18075 -100
rect 18115 -110 18162 15
rect 18210 -35 18258 90
rect 18295 80 18370 90
rect 18295 25 18305 80
rect 18360 25 18370 80
rect 18295 15 18370 25
rect 18195 -45 18270 -35
rect 18195 -100 18205 -45
rect 18260 -100 18270 -45
rect 18195 -110 18270 -100
rect 18308 -110 18355 15
rect 18404 -35 18450 90
rect 18485 80 18560 90
rect 18485 25 18495 80
rect 18550 25 18560 80
rect 18485 15 18560 25
rect 18385 -45 18460 -35
rect 18385 -100 18395 -45
rect 18450 -100 18460 -45
rect 18385 -110 18460 -100
rect 18500 -110 18546 15
rect 18595 -35 18642 90
rect 18675 80 18750 90
rect 18675 25 18685 80
rect 18740 25 18750 80
rect 18675 15 18750 25
rect 18580 -45 18655 -35
rect 18580 -100 18590 -45
rect 18645 -100 18655 -45
rect 18580 -110 18655 -100
rect 18690 -110 18738 15
rect 18788 -35 18835 90
rect 18870 80 18945 90
rect 18870 25 18880 80
rect 18935 25 18945 80
rect 18870 15 18945 25
rect 18770 -45 18845 -35
rect 18770 -100 18780 -45
rect 18835 -100 18845 -45
rect 18770 -110 18845 -100
rect 18884 -110 18930 15
rect 18980 -35 19026 90
rect 19060 80 19135 90
rect 19060 25 19070 80
rect 19125 25 19135 80
rect 19060 15 19135 25
rect 18965 -45 19040 -35
rect 18965 -100 18975 -45
rect 19030 -100 19040 -45
rect 18965 -110 19040 -100
rect 19075 -110 19122 15
rect 19170 -35 19218 90
rect 19255 80 19330 90
rect 19255 25 19265 80
rect 19320 25 19330 80
rect 19255 15 19330 25
rect 19155 -45 19230 -35
rect 19155 -100 19165 -45
rect 19220 -100 19230 -45
rect 19155 -110 19230 -100
rect 19268 -110 19315 15
rect 19364 -35 19410 90
rect 19445 80 19520 90
rect 19445 25 19455 80
rect 19510 25 19520 80
rect 19445 15 19520 25
rect 19350 -45 19425 -35
rect 19350 -100 19360 -45
rect 19415 -100 19425 -45
rect 19350 -110 19425 -100
rect 19460 -110 19506 15
rect 19555 -35 19602 90
rect 19635 80 19710 90
rect 19635 25 19645 80
rect 19700 25 19710 80
rect 19635 15 19710 25
rect 19540 -45 19615 -35
rect 19540 -100 19550 -45
rect 19605 -100 19615 -45
rect 19540 -110 19615 -100
rect 19650 -110 19698 15
rect 19748 -35 19795 90
rect 19830 80 19905 90
rect 19830 25 19840 80
rect 19895 25 19905 80
rect 19830 15 19905 25
rect 19735 -45 19810 -35
rect 19735 -100 19745 -45
rect 19800 -100 19810 -45
rect 19735 -110 19810 -100
rect 19844 -110 19890 15
rect 19940 -35 19986 90
rect 20020 80 20095 90
rect 20020 25 20030 80
rect 20085 25 20095 80
rect 20020 15 20095 25
rect 19925 -45 20000 -35
rect 19925 -100 19935 -45
rect 19990 -100 20000 -45
rect 19925 -110 20000 -100
rect 20035 -110 20082 15
rect 20132 -35 20180 90
rect 20215 80 20290 90
rect 20215 25 20225 80
rect 20280 25 20290 80
rect 20215 15 20290 25
rect 20115 -45 20190 -35
rect 20115 -100 20125 -45
rect 20180 -100 20190 -45
rect 20115 -110 20190 -100
rect 20228 -110 20275 15
rect 20324 -35 20370 90
rect 20405 80 20480 90
rect 20405 25 20415 80
rect 20470 25 20480 80
rect 20405 15 20480 25
rect 20310 -45 20385 -35
rect 20310 -100 20320 -45
rect 20375 -100 20385 -45
rect 20310 -110 20385 -100
rect 20420 -110 20466 15
rect 20515 -35 20562 90
rect 20600 80 20675 90
rect 20600 25 20610 80
rect 20665 25 20675 80
rect 20600 15 20675 25
rect 20500 -45 20575 -35
rect 20500 -100 20510 -45
rect 20565 -100 20575 -45
rect 20500 -110 20575 -100
rect 20610 -110 20658 15
rect 20708 -35 20755 90
rect 20790 80 20865 90
rect 20790 25 20800 80
rect 20855 25 20865 80
rect 20790 15 20865 25
rect 20695 -45 20770 -35
rect 20695 -100 20705 -45
rect 20760 -100 20770 -45
rect 20695 -110 20770 -100
rect 20804 -110 20850 15
rect 20900 -35 20946 90
rect 20980 80 21055 90
rect 20980 25 20990 80
rect 21045 25 21055 80
rect 20980 15 21055 25
rect 20885 -45 20960 -35
rect 20885 -100 20895 -45
rect 20950 -100 20960 -45
rect 20885 -110 20960 -100
rect 20995 -110 21042 15
rect 21090 -35 21138 90
rect 21175 80 21250 90
rect 21175 25 21185 80
rect 21240 25 21250 80
rect 21175 15 21250 25
rect 21075 -45 21150 -35
rect 21075 -100 21085 -45
rect 21140 -100 21150 -45
rect 21075 -110 21150 -100
rect 21188 -110 21235 15
rect 21284 -35 21330 90
rect 21365 80 21440 90
rect 21365 25 21375 80
rect 21430 25 21440 80
rect 21365 15 21440 25
rect 21270 -45 21345 -35
rect 21270 -100 21280 -45
rect 21335 -100 21345 -45
rect 21270 -110 21345 -100
rect 21380 -110 21426 15
rect 21475 -35 21522 90
rect 21555 80 21630 90
rect 21555 25 21565 80
rect 21620 25 21630 80
rect 21555 15 21630 25
rect 21460 -45 21535 -35
rect 21460 -100 21470 -45
rect 21525 -100 21535 -45
rect 21460 -110 21535 -100
rect 21570 -110 21618 15
rect 21668 -35 21715 90
rect 21750 80 21825 90
rect 21750 25 21760 80
rect 21815 25 21825 80
rect 21750 15 21825 25
rect 21650 -45 21725 -35
rect 21650 -100 21660 -45
rect 21715 -100 21725 -45
rect 21650 -110 21725 -100
rect 21764 -110 21810 15
rect 13842 -145 13900 -142
rect 14034 -145 14092 -142
rect 14226 -145 14284 -142
rect 14418 -145 14476 -142
rect 14610 -145 14668 -142
rect 14802 -145 14860 -142
rect 14994 -145 15052 -142
rect 15186 -145 15244 -142
rect 15378 -145 15436 -142
rect 15570 -145 15628 -142
rect 13515 -155 15675 -145
rect 13515 -210 13525 -155
rect 13580 -195 15675 -155
rect 15855 -190 21775 -140
rect 13580 -210 13590 -195
rect 13515 -220 13590 -210
rect 15855 -1840 15905 -190
rect 17435 -565 17870 -530
rect 17435 -1655 17460 -565
rect 17845 -1655 17870 -565
rect 17435 -1675 17870 -1655
<< via1 >>
rect 10210 1190 10605 1720
rect 12170 1185 12575 1720
rect 13740 1190 14120 2280
rect 17455 1190 17840 2280
rect 13525 795 13580 850
rect 9955 685 10010 740
rect 9860 560 9915 615
rect 10150 685 10205 740
rect 10050 560 10105 615
rect 10340 685 10395 740
rect 10240 560 10295 615
rect 10530 685 10585 740
rect 10430 560 10485 615
rect 10720 685 10775 740
rect 10630 560 10685 615
rect 10910 685 10965 740
rect 10820 560 10875 615
rect 11105 685 11160 740
rect 11015 560 11070 615
rect 11300 685 11355 740
rect 11205 560 11260 615
rect 11490 685 11545 740
rect 11395 560 11450 615
rect 11685 685 11740 740
rect 11590 560 11645 615
rect 11780 560 11835 615
rect 12255 685 12310 740
rect 12160 560 12215 615
rect 12445 685 12500 740
rect 12350 560 12405 615
rect 12545 560 12600 615
rect 13795 685 13850 740
rect 13700 560 13755 615
rect 13985 685 14040 740
rect 13890 560 13945 615
rect 14180 685 14235 740
rect 14085 560 14140 615
rect 14370 685 14425 740
rect 14275 560 14330 615
rect 14560 685 14615 740
rect 14470 560 14525 615
rect 14755 685 14810 740
rect 14655 560 14710 615
rect 14945 685 15000 740
rect 14850 560 14905 615
rect 15140 685 15195 740
rect 15040 560 15095 615
rect 15330 685 15385 740
rect 15235 560 15290 615
rect 15520 685 15575 740
rect 15425 560 15480 615
rect 15620 560 15675 615
rect 16095 685 16150 740
rect 15995 560 16050 615
rect 16285 685 16340 740
rect 16185 560 16240 615
rect 16480 685 16535 740
rect 16380 560 16435 615
rect 16670 685 16725 740
rect 16575 560 16630 615
rect 16865 685 16920 740
rect 16765 560 16820 615
rect 17050 685 17105 740
rect 16960 560 17015 615
rect 17250 685 17305 740
rect 17150 560 17205 615
rect 17435 685 17490 740
rect 17345 560 17400 615
rect 17630 685 17685 740
rect 17535 560 17590 615
rect 17825 685 17880 740
rect 17725 560 17780 615
rect 18010 685 18065 740
rect 17920 560 17975 615
rect 18205 685 18260 740
rect 18110 560 18165 615
rect 18395 685 18450 740
rect 18305 560 18360 615
rect 18590 685 18645 740
rect 18495 560 18550 615
rect 18780 685 18835 740
rect 18685 560 18740 615
rect 18975 685 19030 740
rect 18880 560 18935 615
rect 19165 685 19220 740
rect 19070 560 19125 615
rect 19360 685 19415 740
rect 19265 560 19320 615
rect 19550 685 19605 740
rect 19455 560 19510 615
rect 19745 685 19800 740
rect 19645 560 19700 615
rect 19935 685 19990 740
rect 19840 560 19895 615
rect 20125 685 20180 740
rect 20030 560 20085 615
rect 20320 685 20375 740
rect 20225 560 20280 615
rect 20510 685 20565 740
rect 20415 560 20470 615
rect 20705 685 20760 740
rect 20610 560 20665 615
rect 20895 685 20950 740
rect 20800 560 20855 615
rect 21085 685 21140 740
rect 20990 560 21045 615
rect 21280 685 21335 740
rect 21185 560 21240 615
rect 21470 685 21525 740
rect 21375 560 21430 615
rect 21660 685 21715 740
rect 21565 560 21620 615
rect 21760 560 21815 615
rect 9860 25 9915 80
rect 10050 25 10105 80
rect 9955 -100 10010 -45
rect 10240 25 10295 80
rect 10150 -100 10205 -45
rect 10430 25 10485 80
rect 10340 -100 10395 -45
rect 10630 25 10685 80
rect 10530 -100 10585 -45
rect 10820 25 10875 80
rect 10720 -100 10775 -45
rect 11015 25 11070 80
rect 10910 -100 10965 -45
rect 11205 25 11260 80
rect 11105 -100 11160 -45
rect 11395 25 11450 80
rect 11300 -100 11355 -45
rect 11590 25 11645 80
rect 11490 -100 11545 -45
rect 11780 25 11835 80
rect 11685 -100 11740 -45
rect 12160 25 12215 80
rect 12350 25 12405 80
rect 12255 -100 12310 -45
rect 12545 25 12600 80
rect 12445 -100 12500 -45
rect 10205 -1080 10600 -550
rect 12160 -1075 12550 -540
rect 13700 25 13755 80
rect 13890 25 13945 80
rect 13795 -100 13850 -45
rect 14085 25 14140 80
rect 13985 -100 14040 -45
rect 14275 25 14330 80
rect 14180 -100 14235 -45
rect 14470 25 14525 80
rect 14370 -100 14425 -45
rect 14655 25 14710 80
rect 14560 -100 14615 -45
rect 14850 25 14905 80
rect 14755 -100 14810 -45
rect 15040 25 15095 80
rect 14945 -100 15000 -45
rect 15235 25 15290 80
rect 15140 -100 15195 -45
rect 15425 25 15480 80
rect 15330 -100 15385 -45
rect 15620 25 15675 80
rect 15520 -100 15575 -45
rect 15995 25 16050 80
rect 16185 25 16240 80
rect 16095 -100 16150 -45
rect 16380 25 16435 80
rect 16285 -100 16340 -45
rect 16575 25 16630 80
rect 16480 -100 16535 -45
rect 16765 25 16820 80
rect 16670 -100 16725 -45
rect 16960 25 17015 80
rect 16865 -100 16920 -45
rect 17150 25 17205 80
rect 17050 -100 17105 -45
rect 17345 25 17400 80
rect 17250 -100 17305 -45
rect 17535 25 17590 80
rect 17435 -100 17490 -45
rect 17725 25 17780 80
rect 17630 -100 17685 -45
rect 17920 25 17975 80
rect 17825 -100 17880 -45
rect 18110 25 18165 80
rect 18010 -100 18065 -45
rect 18305 25 18360 80
rect 18205 -100 18260 -45
rect 18495 25 18550 80
rect 18395 -100 18450 -45
rect 18685 25 18740 80
rect 18590 -100 18645 -45
rect 18880 25 18935 80
rect 18780 -100 18835 -45
rect 19070 25 19125 80
rect 18975 -100 19030 -45
rect 19265 25 19320 80
rect 19165 -100 19220 -45
rect 19455 25 19510 80
rect 19360 -100 19415 -45
rect 19645 25 19700 80
rect 19550 -100 19605 -45
rect 19840 25 19895 80
rect 19745 -100 19800 -45
rect 20030 25 20085 80
rect 19935 -100 19990 -45
rect 20225 25 20280 80
rect 20125 -100 20180 -45
rect 20415 25 20470 80
rect 20320 -100 20375 -45
rect 20610 25 20665 80
rect 20510 -100 20565 -45
rect 20800 25 20855 80
rect 20705 -100 20760 -45
rect 20990 25 21045 80
rect 20895 -100 20950 -45
rect 21185 25 21240 80
rect 21085 -100 21140 -45
rect 21375 25 21430 80
rect 21280 -100 21335 -45
rect 21565 25 21620 80
rect 21470 -100 21525 -45
rect 21760 25 21815 80
rect 21660 -100 21715 -45
rect 13525 -210 13580 -155
rect 13750 -1655 14135 -560
rect 17460 -1655 17845 -565
<< metal2 >>
rect 13715 2280 14160 2315
rect 10195 1720 10620 1735
rect 10195 1190 10210 1720
rect 10605 1190 10620 1720
rect 10195 1165 10620 1190
rect 12155 1720 12590 1735
rect 12155 1185 12170 1720
rect 12575 1185 12590 1720
rect 12155 1070 12590 1185
rect 13715 1190 13740 2280
rect 14120 1190 14160 2280
rect 13715 1165 14160 1190
rect 17435 2280 17870 2310
rect 17435 1190 17455 2280
rect 17840 1190 17870 2280
rect 17435 1165 17870 1190
rect 12155 1000 13585 1070
rect 8845 975 9985 980
rect 8845 740 11835 975
rect 8845 685 9955 740
rect 10010 685 10150 740
rect 10205 685 10340 740
rect 10395 685 10530 740
rect 10585 685 10720 740
rect 10775 685 10910 740
rect 10965 685 11105 740
rect 11160 685 11300 740
rect 11355 685 11490 740
rect 11545 685 11685 740
rect 11740 685 11835 740
rect 8845 680 11835 685
rect 12155 740 12590 1000
rect 13515 860 13585 1000
rect 13515 850 13590 860
rect 13515 795 13525 850
rect 13580 795 13590 850
rect 13515 785 13590 795
rect 12155 685 12255 740
rect 12310 685 12445 740
rect 12500 685 12590 740
rect 8845 -40 9445 680
rect 12155 675 12590 685
rect 13785 765 13860 775
rect 13785 685 13795 765
rect 13855 695 13860 765
rect 13850 685 13860 695
rect 13785 675 13860 685
rect 13975 765 14050 775
rect 13975 685 13985 765
rect 14045 695 14050 765
rect 14040 685 14050 695
rect 13975 675 14050 685
rect 14170 765 14245 775
rect 14170 685 14180 765
rect 14240 695 14245 765
rect 14235 685 14245 695
rect 14170 675 14245 685
rect 14360 765 14435 775
rect 14360 685 14370 765
rect 14430 695 14435 765
rect 14425 685 14435 695
rect 14360 675 14435 685
rect 14550 765 14625 775
rect 14550 685 14560 765
rect 14620 695 14625 765
rect 14615 685 14625 695
rect 14550 675 14625 685
rect 14745 765 14820 775
rect 14745 685 14755 765
rect 14815 695 14820 765
rect 14810 685 14820 695
rect 14745 675 14820 685
rect 14935 765 15010 775
rect 14935 685 14945 765
rect 15005 695 15010 765
rect 15000 685 15010 695
rect 14935 675 15010 685
rect 15130 765 15205 775
rect 15130 685 15140 765
rect 15200 695 15205 765
rect 15195 685 15205 695
rect 15130 675 15205 685
rect 15320 765 15395 775
rect 15320 685 15330 765
rect 15390 695 15395 765
rect 15385 685 15395 695
rect 15320 675 15395 685
rect 15510 765 15585 775
rect 15510 685 15520 765
rect 15580 695 15585 765
rect 15575 685 15585 695
rect 15510 675 15585 685
rect 16085 765 16160 775
rect 16085 695 16090 765
rect 16085 685 16095 695
rect 16150 685 16160 765
rect 16085 675 16160 685
rect 16275 765 16350 775
rect 16275 695 16280 765
rect 16275 685 16285 695
rect 16340 685 16350 765
rect 16275 675 16350 685
rect 16470 765 16545 775
rect 16470 695 16475 765
rect 16470 685 16480 695
rect 16535 685 16545 765
rect 16470 675 16545 685
rect 16660 765 16735 775
rect 16660 695 16665 765
rect 16660 685 16670 695
rect 16725 685 16735 765
rect 16660 675 16735 685
rect 16855 765 16930 775
rect 16855 695 16860 765
rect 16855 685 16865 695
rect 16920 685 16930 765
rect 16855 675 16930 685
rect 17040 765 17115 775
rect 17040 695 17045 765
rect 17040 685 17050 695
rect 17105 685 17115 765
rect 17040 675 17115 685
rect 17240 765 17315 775
rect 17240 695 17245 765
rect 17240 685 17250 695
rect 17305 685 17315 765
rect 17240 675 17315 685
rect 17425 765 17500 775
rect 17425 695 17430 765
rect 17425 685 17435 695
rect 17490 685 17500 765
rect 17425 675 17500 685
rect 17620 765 17695 775
rect 17620 695 17625 765
rect 17620 685 17630 695
rect 17685 685 17695 765
rect 17620 675 17695 685
rect 17815 765 17890 775
rect 17815 695 17820 765
rect 17815 685 17825 695
rect 17880 685 17890 765
rect 17815 675 17890 685
rect 18000 765 18075 775
rect 18000 695 18005 765
rect 18000 685 18010 695
rect 18065 685 18075 765
rect 18000 675 18075 685
rect 18195 765 18270 775
rect 18195 695 18200 765
rect 18195 685 18205 695
rect 18260 685 18270 765
rect 18195 675 18270 685
rect 18385 765 18460 775
rect 18385 695 18390 765
rect 18385 685 18395 695
rect 18450 685 18460 765
rect 18385 675 18460 685
rect 18580 765 18655 775
rect 18580 695 18585 765
rect 18580 685 18590 695
rect 18645 685 18655 765
rect 18580 675 18655 685
rect 18770 765 18845 775
rect 18770 695 18775 765
rect 18770 685 18780 695
rect 18835 685 18845 765
rect 18770 675 18845 685
rect 18965 765 19040 775
rect 18965 695 18970 765
rect 18965 685 18975 695
rect 19030 685 19040 765
rect 18965 675 19040 685
rect 19155 765 19230 775
rect 19155 695 19160 765
rect 19155 685 19165 695
rect 19220 685 19230 765
rect 19155 675 19230 685
rect 19350 765 19425 775
rect 19350 695 19355 765
rect 19350 685 19360 695
rect 19415 685 19425 765
rect 19350 675 19425 685
rect 19540 765 19615 775
rect 19540 695 19545 765
rect 19540 685 19550 695
rect 19605 685 19615 765
rect 19540 675 19615 685
rect 19735 765 19810 775
rect 19735 695 19740 765
rect 19735 685 19745 695
rect 19800 685 19810 765
rect 19735 675 19810 685
rect 19925 765 20000 775
rect 19925 695 19930 765
rect 19925 685 19935 695
rect 19990 685 20000 765
rect 19925 675 20000 685
rect 20115 765 20190 775
rect 20115 695 20120 765
rect 20115 685 20125 695
rect 20180 685 20190 765
rect 20115 675 20190 685
rect 20310 765 20385 775
rect 20310 695 20315 765
rect 20310 685 20320 695
rect 20375 685 20385 765
rect 20310 675 20385 685
rect 20500 765 20575 775
rect 20500 695 20505 765
rect 20500 685 20510 695
rect 20565 685 20575 765
rect 20500 675 20575 685
rect 20695 765 20770 775
rect 20695 695 20700 765
rect 20695 685 20705 695
rect 20760 685 20770 765
rect 20695 675 20770 685
rect 20885 765 20960 775
rect 20885 695 20890 765
rect 20885 685 20895 695
rect 20950 685 20960 765
rect 20885 675 20960 685
rect 21075 765 21150 775
rect 21075 695 21080 765
rect 21075 685 21085 695
rect 21140 685 21150 765
rect 21075 675 21150 685
rect 21270 765 21345 775
rect 21270 695 21275 765
rect 21270 685 21280 695
rect 21335 685 21345 765
rect 21270 675 21345 685
rect 21460 765 21535 775
rect 21460 695 21465 765
rect 21460 685 21470 695
rect 21525 685 21535 765
rect 21460 675 21535 685
rect 21650 765 21725 775
rect 21650 695 21655 765
rect 21650 685 21660 695
rect 21715 685 21725 765
rect 21650 675 21725 685
rect 12150 620 12225 625
rect 12340 620 12415 625
rect 12535 620 12610 625
rect 9850 615 12610 620
rect 9850 560 9860 615
rect 9915 560 10050 615
rect 10105 560 10240 615
rect 10295 560 10430 615
rect 10485 560 10630 615
rect 10685 560 10820 615
rect 10875 560 11015 615
rect 11070 560 11205 615
rect 11260 560 11395 615
rect 11450 560 11590 615
rect 11645 560 11780 615
rect 11835 560 12160 615
rect 12215 560 12350 615
rect 12405 560 12545 615
rect 12600 560 12610 615
rect 9850 80 12610 560
rect 13690 615 13765 625
rect 13690 535 13700 615
rect 13755 605 13765 615
rect 13760 535 13765 605
rect 13690 525 13765 535
rect 13880 615 13955 625
rect 13880 535 13890 615
rect 13945 605 13955 615
rect 13950 535 13955 605
rect 13880 525 13955 535
rect 14075 615 14150 625
rect 14075 535 14085 615
rect 14140 605 14150 615
rect 14145 535 14150 605
rect 14075 525 14150 535
rect 14265 615 14340 625
rect 14265 535 14275 615
rect 14330 605 14340 615
rect 14335 535 14340 605
rect 14265 525 14340 535
rect 14460 615 14535 625
rect 14460 535 14470 615
rect 14525 605 14535 615
rect 14530 535 14535 605
rect 14460 525 14535 535
rect 14645 615 14720 625
rect 14645 535 14655 615
rect 14710 605 14720 615
rect 14715 535 14720 605
rect 14645 525 14720 535
rect 14840 615 14915 625
rect 14840 535 14850 615
rect 14905 605 14915 615
rect 14910 535 14915 605
rect 14840 525 14915 535
rect 15030 615 15105 625
rect 15030 535 15040 615
rect 15095 605 15105 615
rect 15100 535 15105 605
rect 15030 525 15105 535
rect 15225 615 15300 625
rect 15225 535 15235 615
rect 15290 605 15300 615
rect 15295 535 15300 605
rect 15225 525 15300 535
rect 15415 615 15490 625
rect 15415 535 15425 615
rect 15480 605 15490 615
rect 15485 535 15490 605
rect 15415 525 15490 535
rect 15610 615 15685 625
rect 15610 535 15620 615
rect 15675 605 15685 615
rect 15680 535 15685 605
rect 15610 525 15685 535
rect 15985 615 16060 625
rect 15985 535 15995 615
rect 16050 605 16060 615
rect 16055 535 16060 605
rect 15985 525 16060 535
rect 16175 615 16250 625
rect 16175 535 16185 615
rect 16240 605 16250 615
rect 16245 535 16250 605
rect 16175 525 16250 535
rect 16370 615 16445 625
rect 16370 535 16380 615
rect 16435 605 16445 615
rect 16440 535 16445 605
rect 16370 525 16445 535
rect 16565 615 16640 625
rect 16565 535 16575 615
rect 16630 605 16640 615
rect 16635 535 16640 605
rect 16565 525 16640 535
rect 16755 615 16830 625
rect 16755 535 16765 615
rect 16820 605 16830 615
rect 16825 535 16830 605
rect 16755 525 16830 535
rect 16950 615 17025 625
rect 16950 535 16960 615
rect 17015 605 17025 615
rect 17020 535 17025 605
rect 16950 525 17025 535
rect 17140 615 17215 625
rect 17140 535 17150 615
rect 17205 605 17215 615
rect 17210 535 17215 605
rect 17140 525 17215 535
rect 17335 615 17410 625
rect 17335 535 17345 615
rect 17400 605 17410 615
rect 17405 535 17410 605
rect 17335 525 17410 535
rect 17525 615 17600 625
rect 17525 535 17535 615
rect 17590 605 17600 615
rect 17595 535 17600 605
rect 17525 525 17600 535
rect 17715 615 17790 625
rect 17715 535 17725 615
rect 17780 605 17790 615
rect 17785 535 17790 605
rect 17715 525 17790 535
rect 17910 615 17985 625
rect 17910 535 17920 615
rect 17975 605 17985 615
rect 17980 535 17985 605
rect 17910 525 17985 535
rect 18100 615 18175 625
rect 18100 535 18110 615
rect 18165 605 18175 615
rect 18170 535 18175 605
rect 18100 525 18175 535
rect 18295 615 18370 625
rect 18295 535 18305 615
rect 18360 605 18370 615
rect 18365 535 18370 605
rect 18295 525 18370 535
rect 18485 615 18560 625
rect 18485 535 18495 615
rect 18550 605 18560 615
rect 18555 535 18560 605
rect 18485 525 18560 535
rect 18675 615 18750 625
rect 18675 535 18685 615
rect 18740 605 18750 615
rect 18745 535 18750 605
rect 18675 525 18750 535
rect 18870 615 18945 625
rect 18870 535 18880 615
rect 18935 605 18945 615
rect 18940 535 18945 605
rect 18870 525 18945 535
rect 19060 615 19135 625
rect 19060 535 19070 615
rect 19125 605 19135 615
rect 19130 535 19135 605
rect 19060 525 19135 535
rect 19255 615 19330 625
rect 19255 535 19265 615
rect 19320 605 19330 615
rect 19325 535 19330 605
rect 19255 525 19330 535
rect 19445 615 19520 625
rect 19445 535 19455 615
rect 19510 605 19520 615
rect 19515 535 19520 605
rect 19445 525 19520 535
rect 19635 615 19710 625
rect 19635 535 19645 615
rect 19700 605 19710 615
rect 19705 535 19710 605
rect 19635 525 19710 535
rect 19830 615 19905 625
rect 19830 535 19840 615
rect 19895 605 19905 615
rect 19900 535 19905 605
rect 19830 525 19905 535
rect 20020 615 20095 625
rect 20020 535 20030 615
rect 20085 605 20095 615
rect 20090 535 20095 605
rect 20020 525 20095 535
rect 20215 615 20290 625
rect 20215 535 20225 615
rect 20280 605 20290 615
rect 20285 535 20290 605
rect 20215 525 20290 535
rect 20405 615 20480 625
rect 20405 535 20415 615
rect 20470 605 20480 615
rect 20475 535 20480 605
rect 20405 525 20480 535
rect 20600 615 20675 625
rect 20600 535 20610 615
rect 20665 605 20675 615
rect 20670 535 20675 605
rect 20600 525 20675 535
rect 20790 615 20865 625
rect 20790 535 20800 615
rect 20855 605 20865 615
rect 20860 535 20865 605
rect 20790 525 20865 535
rect 20980 615 21055 625
rect 20980 535 20990 615
rect 21045 605 21055 615
rect 21050 535 21055 605
rect 20980 525 21055 535
rect 21175 615 21250 625
rect 21175 535 21185 615
rect 21240 605 21250 615
rect 21245 535 21250 605
rect 21175 525 21250 535
rect 21365 615 21440 625
rect 21365 535 21375 615
rect 21430 605 21440 615
rect 21435 535 21440 605
rect 21365 525 21440 535
rect 21555 615 21630 625
rect 21555 535 21565 615
rect 21620 605 21630 615
rect 21625 535 21630 605
rect 21555 525 21630 535
rect 21750 615 21825 625
rect 21750 535 21760 615
rect 21815 605 21825 615
rect 21820 535 21825 605
rect 21750 525 21825 535
rect 9850 25 9860 80
rect 9915 25 10050 80
rect 10105 25 10240 80
rect 10295 25 10430 80
rect 10485 25 10630 80
rect 10685 25 10820 80
rect 10875 25 11015 80
rect 11070 25 11205 80
rect 11260 25 11395 80
rect 11450 25 11590 80
rect 11645 25 11780 80
rect 11835 25 12160 80
rect 12215 25 12350 80
rect 12405 25 12545 80
rect 12600 25 12610 80
rect 9850 20 12610 25
rect 12150 15 12225 20
rect 12340 15 12415 20
rect 12535 15 12610 20
rect 13690 105 13765 115
rect 13690 25 13700 105
rect 13760 35 13765 105
rect 13755 25 13765 35
rect 13690 15 13765 25
rect 13880 105 13955 115
rect 13880 25 13890 105
rect 13950 35 13955 105
rect 13945 25 13955 35
rect 13880 15 13955 25
rect 14075 105 14150 115
rect 14075 25 14085 105
rect 14145 35 14150 105
rect 14140 25 14150 35
rect 14075 15 14150 25
rect 14265 105 14340 115
rect 14265 25 14275 105
rect 14335 35 14340 105
rect 14330 25 14340 35
rect 14265 15 14340 25
rect 14460 105 14535 115
rect 14460 25 14470 105
rect 14530 35 14535 105
rect 14525 25 14535 35
rect 14460 15 14535 25
rect 14645 105 14720 115
rect 14645 25 14655 105
rect 14715 35 14720 105
rect 14710 25 14720 35
rect 14645 15 14720 25
rect 14840 105 14915 115
rect 14840 25 14850 105
rect 14910 35 14915 105
rect 14905 25 14915 35
rect 14840 15 14915 25
rect 15030 105 15105 115
rect 15030 25 15040 105
rect 15100 35 15105 105
rect 15095 25 15105 35
rect 15030 15 15105 25
rect 15225 105 15300 115
rect 15225 25 15235 105
rect 15295 35 15300 105
rect 15290 25 15300 35
rect 15225 15 15300 25
rect 15415 105 15490 115
rect 15415 25 15425 105
rect 15485 35 15490 105
rect 15480 25 15490 35
rect 15415 15 15490 25
rect 15610 105 15685 115
rect 15610 25 15620 105
rect 15680 35 15685 105
rect 15675 25 15685 35
rect 15610 15 15685 25
rect 15985 105 16060 115
rect 15985 25 15995 105
rect 16055 35 16060 105
rect 16050 25 16060 35
rect 15985 15 16060 25
rect 16175 105 16250 115
rect 16175 25 16185 105
rect 16245 35 16250 105
rect 16240 25 16250 35
rect 16175 15 16250 25
rect 16370 105 16445 115
rect 16370 25 16380 105
rect 16440 35 16445 105
rect 16435 25 16445 35
rect 16370 15 16445 25
rect 16565 105 16640 115
rect 16565 25 16575 105
rect 16635 35 16640 105
rect 16630 25 16640 35
rect 16565 15 16640 25
rect 16755 105 16830 115
rect 16755 25 16765 105
rect 16825 35 16830 105
rect 16820 25 16830 35
rect 16755 15 16830 25
rect 16950 105 17025 115
rect 16950 25 16960 105
rect 17020 35 17025 105
rect 17015 25 17025 35
rect 16950 15 17025 25
rect 17140 105 17215 115
rect 17140 25 17150 105
rect 17210 35 17215 105
rect 17205 25 17215 35
rect 17140 15 17215 25
rect 17335 105 17410 115
rect 17335 25 17345 105
rect 17405 35 17410 105
rect 17400 25 17410 35
rect 17335 15 17410 25
rect 17525 105 17600 115
rect 17525 25 17535 105
rect 17595 35 17600 105
rect 17590 25 17600 35
rect 17525 15 17600 25
rect 17715 105 17790 115
rect 17715 25 17725 105
rect 17785 35 17790 105
rect 17780 25 17790 35
rect 17715 15 17790 25
rect 17910 105 17985 115
rect 17910 25 17920 105
rect 17980 35 17985 105
rect 17975 25 17985 35
rect 17910 15 17985 25
rect 18100 105 18175 115
rect 18100 25 18110 105
rect 18170 35 18175 105
rect 18165 25 18175 35
rect 18100 15 18175 25
rect 18295 105 18370 115
rect 18295 25 18305 105
rect 18365 35 18370 105
rect 18360 25 18370 35
rect 18295 15 18370 25
rect 18485 105 18560 115
rect 18485 25 18495 105
rect 18555 35 18560 105
rect 18550 25 18560 35
rect 18485 15 18560 25
rect 18675 105 18750 115
rect 18675 25 18685 105
rect 18745 35 18750 105
rect 18740 25 18750 35
rect 18675 15 18750 25
rect 18870 105 18945 115
rect 18870 25 18880 105
rect 18940 35 18945 105
rect 18935 25 18945 35
rect 18870 15 18945 25
rect 19060 105 19135 115
rect 19060 25 19070 105
rect 19130 35 19135 105
rect 19125 25 19135 35
rect 19060 15 19135 25
rect 19255 105 19330 115
rect 19255 25 19265 105
rect 19325 35 19330 105
rect 19320 25 19330 35
rect 19255 15 19330 25
rect 19445 105 19520 115
rect 19445 25 19455 105
rect 19515 35 19520 105
rect 19510 25 19520 35
rect 19445 15 19520 25
rect 19635 105 19710 115
rect 19635 25 19645 105
rect 19705 35 19710 105
rect 19700 25 19710 35
rect 19635 15 19710 25
rect 19830 105 19905 115
rect 19830 25 19840 105
rect 19900 35 19905 105
rect 19895 25 19905 35
rect 19830 15 19905 25
rect 20020 105 20095 115
rect 20020 25 20030 105
rect 20090 35 20095 105
rect 20085 25 20095 35
rect 20020 15 20095 25
rect 20215 105 20290 115
rect 20215 25 20225 105
rect 20285 35 20290 105
rect 20280 25 20290 35
rect 20215 15 20290 25
rect 20405 105 20480 115
rect 20405 25 20415 105
rect 20475 35 20480 105
rect 20470 25 20480 35
rect 20405 15 20480 25
rect 20600 105 20675 115
rect 20600 25 20610 105
rect 20670 35 20675 105
rect 20665 25 20675 35
rect 20600 15 20675 25
rect 20790 105 20865 115
rect 20790 25 20800 105
rect 20860 35 20865 105
rect 20855 25 20865 35
rect 20790 15 20865 25
rect 20980 105 21055 115
rect 20980 25 20990 105
rect 21050 35 21055 105
rect 21045 25 21055 35
rect 20980 15 21055 25
rect 21175 105 21250 115
rect 21175 25 21185 105
rect 21245 35 21250 105
rect 21240 25 21250 35
rect 21175 15 21250 25
rect 21365 105 21440 115
rect 21365 25 21375 105
rect 21435 35 21440 105
rect 21430 25 21440 35
rect 21365 15 21440 25
rect 21555 105 21630 115
rect 21555 25 21565 105
rect 21625 35 21630 105
rect 21620 25 21630 35
rect 21555 15 21630 25
rect 21750 105 21825 115
rect 21750 25 21760 105
rect 21820 35 21825 105
rect 21815 25 21825 35
rect 21750 15 21825 25
rect 8845 -45 11835 -40
rect 8845 -100 9955 -45
rect 10010 -100 10150 -45
rect 10205 -100 10340 -45
rect 10395 -100 10530 -45
rect 10585 -100 10720 -45
rect 10775 -100 10910 -45
rect 10965 -100 11105 -45
rect 11160 -100 11300 -45
rect 11355 -100 11490 -45
rect 11545 -100 11685 -45
rect 11740 -100 11835 -45
rect 8845 -340 11835 -100
rect 12140 -45 12565 -35
rect 12140 -100 12255 -45
rect 12310 -100 12445 -45
rect 12500 -100 12565 -45
rect 8845 -1300 9445 -340
rect 12140 -370 12565 -100
rect 13785 -45 13860 -35
rect 13785 -125 13795 -45
rect 13850 -55 13860 -45
rect 13855 -125 13860 -55
rect 13785 -135 13860 -125
rect 13975 -45 14050 -35
rect 13975 -125 13985 -45
rect 14040 -55 14050 -45
rect 14045 -125 14050 -55
rect 13975 -135 14050 -125
rect 14170 -45 14245 -35
rect 14170 -125 14180 -45
rect 14235 -55 14245 -45
rect 14240 -125 14245 -55
rect 14170 -135 14245 -125
rect 14360 -45 14435 -35
rect 14360 -125 14370 -45
rect 14425 -55 14435 -45
rect 14430 -125 14435 -55
rect 14360 -135 14435 -125
rect 14550 -45 14625 -35
rect 14550 -125 14560 -45
rect 14615 -55 14625 -45
rect 14620 -125 14625 -55
rect 14550 -135 14625 -125
rect 14745 -45 14820 -35
rect 14745 -125 14755 -45
rect 14810 -55 14820 -45
rect 14815 -125 14820 -55
rect 14745 -135 14820 -125
rect 14935 -45 15010 -35
rect 14935 -125 14945 -45
rect 15000 -55 15010 -45
rect 15005 -125 15010 -55
rect 14935 -135 15010 -125
rect 15130 -45 15205 -35
rect 15130 -125 15140 -45
rect 15195 -55 15205 -45
rect 15200 -125 15205 -55
rect 15130 -135 15205 -125
rect 15320 -45 15395 -35
rect 15320 -125 15330 -45
rect 15385 -55 15395 -45
rect 15390 -125 15395 -55
rect 15320 -135 15395 -125
rect 15510 -45 15585 -35
rect 15510 -125 15520 -45
rect 15575 -55 15585 -45
rect 15580 -125 15585 -55
rect 15510 -135 15585 -125
rect 16085 -45 16160 -35
rect 16085 -55 16095 -45
rect 16085 -125 16090 -55
rect 16150 -125 16160 -45
rect 16085 -135 16160 -125
rect 16275 -45 16350 -35
rect 16275 -55 16285 -45
rect 16275 -125 16280 -55
rect 16340 -125 16350 -45
rect 16275 -135 16350 -125
rect 16470 -45 16545 -35
rect 16470 -55 16480 -45
rect 16470 -125 16475 -55
rect 16535 -125 16545 -45
rect 16470 -135 16545 -125
rect 16660 -45 16735 -35
rect 16660 -55 16670 -45
rect 16660 -125 16665 -55
rect 16725 -125 16735 -45
rect 16660 -135 16735 -125
rect 16855 -45 16930 -35
rect 16855 -55 16865 -45
rect 16855 -125 16860 -55
rect 16920 -125 16930 -45
rect 16855 -135 16930 -125
rect 17040 -45 17115 -35
rect 17040 -55 17050 -45
rect 17040 -125 17045 -55
rect 17105 -125 17115 -45
rect 17040 -135 17115 -125
rect 17240 -45 17315 -35
rect 17240 -55 17250 -45
rect 17240 -125 17245 -55
rect 17305 -125 17315 -45
rect 17240 -135 17315 -125
rect 17425 -45 17500 -35
rect 17425 -55 17435 -45
rect 17425 -125 17430 -55
rect 17490 -125 17500 -45
rect 17425 -135 17500 -125
rect 17620 -45 17695 -35
rect 17620 -55 17630 -45
rect 17620 -125 17625 -55
rect 17685 -125 17695 -45
rect 17620 -135 17695 -125
rect 17815 -45 17890 -35
rect 17815 -55 17825 -45
rect 17815 -125 17820 -55
rect 17880 -125 17890 -45
rect 17815 -135 17890 -125
rect 18000 -45 18075 -35
rect 18000 -55 18010 -45
rect 18000 -125 18005 -55
rect 18065 -125 18075 -45
rect 18000 -135 18075 -125
rect 18195 -45 18270 -35
rect 18195 -55 18205 -45
rect 18195 -125 18200 -55
rect 18260 -125 18270 -45
rect 18195 -135 18270 -125
rect 18385 -45 18460 -35
rect 18385 -55 18395 -45
rect 18385 -125 18390 -55
rect 18450 -125 18460 -45
rect 18385 -135 18460 -125
rect 18580 -45 18655 -35
rect 18580 -55 18590 -45
rect 18580 -125 18585 -55
rect 18645 -125 18655 -45
rect 18580 -135 18655 -125
rect 18770 -45 18845 -35
rect 18770 -55 18780 -45
rect 18770 -125 18775 -55
rect 18835 -125 18845 -45
rect 18770 -135 18845 -125
rect 18965 -45 19040 -35
rect 18965 -55 18975 -45
rect 18965 -125 18970 -55
rect 19030 -125 19040 -45
rect 18965 -135 19040 -125
rect 19155 -45 19230 -35
rect 19155 -55 19165 -45
rect 19155 -125 19160 -55
rect 19220 -125 19230 -45
rect 19155 -135 19230 -125
rect 19350 -45 19425 -35
rect 19350 -55 19360 -45
rect 19350 -125 19355 -55
rect 19415 -125 19425 -45
rect 19350 -135 19425 -125
rect 19540 -45 19615 -35
rect 19540 -55 19550 -45
rect 19540 -125 19545 -55
rect 19605 -125 19615 -45
rect 19540 -135 19615 -125
rect 19735 -45 19810 -35
rect 19735 -55 19745 -45
rect 19735 -125 19740 -55
rect 19800 -125 19810 -45
rect 19735 -135 19810 -125
rect 19925 -45 20000 -35
rect 19925 -55 19935 -45
rect 19925 -125 19930 -55
rect 19990 -125 20000 -45
rect 19925 -135 20000 -125
rect 20115 -45 20190 -35
rect 20115 -55 20125 -45
rect 20115 -125 20120 -55
rect 20180 -125 20190 -45
rect 20115 -135 20190 -125
rect 20310 -45 20385 -35
rect 20310 -55 20320 -45
rect 20310 -125 20315 -55
rect 20375 -125 20385 -45
rect 20310 -135 20385 -125
rect 20500 -45 20575 -35
rect 20500 -55 20510 -45
rect 20500 -125 20505 -55
rect 20565 -125 20575 -45
rect 20500 -135 20575 -125
rect 20695 -45 20770 -35
rect 20695 -55 20705 -45
rect 20695 -125 20700 -55
rect 20760 -125 20770 -45
rect 20695 -135 20770 -125
rect 20885 -45 20960 -35
rect 20885 -55 20895 -45
rect 20885 -125 20890 -55
rect 20950 -125 20960 -45
rect 20885 -135 20960 -125
rect 21075 -45 21150 -35
rect 21075 -55 21085 -45
rect 21075 -125 21080 -55
rect 21140 -125 21150 -45
rect 21075 -135 21150 -125
rect 21270 -45 21345 -35
rect 21270 -55 21280 -45
rect 21270 -125 21275 -55
rect 21335 -125 21345 -45
rect 21270 -135 21345 -125
rect 21460 -45 21535 -35
rect 21460 -55 21470 -45
rect 21460 -125 21465 -55
rect 21525 -125 21535 -45
rect 21460 -135 21535 -125
rect 21650 -45 21725 -35
rect 21650 -55 21660 -45
rect 21650 -125 21655 -55
rect 21715 -125 21725 -45
rect 21650 -135 21725 -125
rect 13515 -155 13590 -145
rect 13515 -210 13525 -155
rect 13580 -210 13590 -155
rect 13515 -370 13590 -210
rect 12140 -440 13590 -370
rect 10190 -550 10615 -520
rect 10190 -1080 10205 -550
rect 10600 -1080 10615 -550
rect 10190 -1090 10615 -1080
rect 12140 -540 12565 -440
rect 12140 -1075 12160 -540
rect 12550 -1075 12565 -540
rect 12140 -1090 12565 -1075
rect 13725 -560 14165 -520
rect 13725 -1655 13750 -560
rect 14135 -1655 14165 -560
rect 13725 -1675 14165 -1655
rect 17435 -565 17870 -530
rect 17435 -1655 17460 -565
rect 17845 -1655 17870 -565
rect 17435 -1675 17870 -1655
<< via2 >>
rect 10210 1190 10605 1720
rect 13740 1190 14120 2280
rect 17455 1190 17840 2280
rect 13795 740 13855 765
rect 13795 695 13850 740
rect 13850 695 13855 740
rect 13985 740 14045 765
rect 13985 695 14040 740
rect 14040 695 14045 740
rect 14180 740 14240 765
rect 14180 695 14235 740
rect 14235 695 14240 740
rect 14370 740 14430 765
rect 14370 695 14425 740
rect 14425 695 14430 740
rect 14560 740 14620 765
rect 14560 695 14615 740
rect 14615 695 14620 740
rect 14755 740 14815 765
rect 14755 695 14810 740
rect 14810 695 14815 740
rect 14945 740 15005 765
rect 14945 695 15000 740
rect 15000 695 15005 740
rect 15140 740 15200 765
rect 15140 695 15195 740
rect 15195 695 15200 740
rect 15330 740 15390 765
rect 15330 695 15385 740
rect 15385 695 15390 740
rect 15520 740 15580 765
rect 15520 695 15575 740
rect 15575 695 15580 740
rect 16090 740 16150 765
rect 16090 695 16095 740
rect 16095 695 16150 740
rect 16280 740 16340 765
rect 16280 695 16285 740
rect 16285 695 16340 740
rect 16475 740 16535 765
rect 16475 695 16480 740
rect 16480 695 16535 740
rect 16665 740 16725 765
rect 16665 695 16670 740
rect 16670 695 16725 740
rect 16860 740 16920 765
rect 16860 695 16865 740
rect 16865 695 16920 740
rect 17045 740 17105 765
rect 17045 695 17050 740
rect 17050 695 17105 740
rect 17245 740 17305 765
rect 17245 695 17250 740
rect 17250 695 17305 740
rect 17430 740 17490 765
rect 17430 695 17435 740
rect 17435 695 17490 740
rect 17625 740 17685 765
rect 17625 695 17630 740
rect 17630 695 17685 740
rect 17820 740 17880 765
rect 17820 695 17825 740
rect 17825 695 17880 740
rect 18005 740 18065 765
rect 18005 695 18010 740
rect 18010 695 18065 740
rect 18200 740 18260 765
rect 18200 695 18205 740
rect 18205 695 18260 740
rect 18390 740 18450 765
rect 18390 695 18395 740
rect 18395 695 18450 740
rect 18585 740 18645 765
rect 18585 695 18590 740
rect 18590 695 18645 740
rect 18775 740 18835 765
rect 18775 695 18780 740
rect 18780 695 18835 740
rect 18970 740 19030 765
rect 18970 695 18975 740
rect 18975 695 19030 740
rect 19160 740 19220 765
rect 19160 695 19165 740
rect 19165 695 19220 740
rect 19355 740 19415 765
rect 19355 695 19360 740
rect 19360 695 19415 740
rect 19545 740 19605 765
rect 19545 695 19550 740
rect 19550 695 19605 740
rect 19740 740 19800 765
rect 19740 695 19745 740
rect 19745 695 19800 740
rect 19930 740 19990 765
rect 19930 695 19935 740
rect 19935 695 19990 740
rect 20120 740 20180 765
rect 20120 695 20125 740
rect 20125 695 20180 740
rect 20315 740 20375 765
rect 20315 695 20320 740
rect 20320 695 20375 740
rect 20505 740 20565 765
rect 20505 695 20510 740
rect 20510 695 20565 740
rect 20700 740 20760 765
rect 20700 695 20705 740
rect 20705 695 20760 740
rect 20890 740 20950 765
rect 20890 695 20895 740
rect 20895 695 20950 740
rect 21080 740 21140 765
rect 21080 695 21085 740
rect 21085 695 21140 740
rect 21275 740 21335 765
rect 21275 695 21280 740
rect 21280 695 21335 740
rect 21465 740 21525 765
rect 21465 695 21470 740
rect 21470 695 21525 740
rect 21655 740 21715 765
rect 21655 695 21660 740
rect 21660 695 21715 740
rect 13700 560 13755 605
rect 13755 560 13760 605
rect 13700 535 13760 560
rect 13890 560 13945 605
rect 13945 560 13950 605
rect 13890 535 13950 560
rect 14085 560 14140 605
rect 14140 560 14145 605
rect 14085 535 14145 560
rect 14275 560 14330 605
rect 14330 560 14335 605
rect 14275 535 14335 560
rect 14470 560 14525 605
rect 14525 560 14530 605
rect 14470 535 14530 560
rect 14655 560 14710 605
rect 14710 560 14715 605
rect 14655 535 14715 560
rect 14850 560 14905 605
rect 14905 560 14910 605
rect 14850 535 14910 560
rect 15040 560 15095 605
rect 15095 560 15100 605
rect 15040 535 15100 560
rect 15235 560 15290 605
rect 15290 560 15295 605
rect 15235 535 15295 560
rect 15425 560 15480 605
rect 15480 560 15485 605
rect 15425 535 15485 560
rect 15620 560 15675 605
rect 15675 560 15680 605
rect 15620 535 15680 560
rect 15995 560 16050 605
rect 16050 560 16055 605
rect 15995 535 16055 560
rect 16185 560 16240 605
rect 16240 560 16245 605
rect 16185 535 16245 560
rect 16380 560 16435 605
rect 16435 560 16440 605
rect 16380 535 16440 560
rect 16575 560 16630 605
rect 16630 560 16635 605
rect 16575 535 16635 560
rect 16765 560 16820 605
rect 16820 560 16825 605
rect 16765 535 16825 560
rect 16960 560 17015 605
rect 17015 560 17020 605
rect 16960 535 17020 560
rect 17150 560 17205 605
rect 17205 560 17210 605
rect 17150 535 17210 560
rect 17345 560 17400 605
rect 17400 560 17405 605
rect 17345 535 17405 560
rect 17535 560 17590 605
rect 17590 560 17595 605
rect 17535 535 17595 560
rect 17725 560 17780 605
rect 17780 560 17785 605
rect 17725 535 17785 560
rect 17920 560 17975 605
rect 17975 560 17980 605
rect 17920 535 17980 560
rect 18110 560 18165 605
rect 18165 560 18170 605
rect 18110 535 18170 560
rect 18305 560 18360 605
rect 18360 560 18365 605
rect 18305 535 18365 560
rect 18495 560 18550 605
rect 18550 560 18555 605
rect 18495 535 18555 560
rect 18685 560 18740 605
rect 18740 560 18745 605
rect 18685 535 18745 560
rect 18880 560 18935 605
rect 18935 560 18940 605
rect 18880 535 18940 560
rect 19070 560 19125 605
rect 19125 560 19130 605
rect 19070 535 19130 560
rect 19265 560 19320 605
rect 19320 560 19325 605
rect 19265 535 19325 560
rect 19455 560 19510 605
rect 19510 560 19515 605
rect 19455 535 19515 560
rect 19645 560 19700 605
rect 19700 560 19705 605
rect 19645 535 19705 560
rect 19840 560 19895 605
rect 19895 560 19900 605
rect 19840 535 19900 560
rect 20030 560 20085 605
rect 20085 560 20090 605
rect 20030 535 20090 560
rect 20225 560 20280 605
rect 20280 560 20285 605
rect 20225 535 20285 560
rect 20415 560 20470 605
rect 20470 560 20475 605
rect 20415 535 20475 560
rect 20610 560 20665 605
rect 20665 560 20670 605
rect 20610 535 20670 560
rect 20800 560 20855 605
rect 20855 560 20860 605
rect 20800 535 20860 560
rect 20990 560 21045 605
rect 21045 560 21050 605
rect 20990 535 21050 560
rect 21185 560 21240 605
rect 21240 560 21245 605
rect 21185 535 21245 560
rect 21375 560 21430 605
rect 21430 560 21435 605
rect 21375 535 21435 560
rect 21565 560 21620 605
rect 21620 560 21625 605
rect 21565 535 21625 560
rect 21760 560 21815 605
rect 21815 560 21820 605
rect 21760 535 21820 560
rect 13700 80 13760 105
rect 13700 35 13755 80
rect 13755 35 13760 80
rect 13890 80 13950 105
rect 13890 35 13945 80
rect 13945 35 13950 80
rect 14085 80 14145 105
rect 14085 35 14140 80
rect 14140 35 14145 80
rect 14275 80 14335 105
rect 14275 35 14330 80
rect 14330 35 14335 80
rect 14470 80 14530 105
rect 14470 35 14525 80
rect 14525 35 14530 80
rect 14655 80 14715 105
rect 14655 35 14710 80
rect 14710 35 14715 80
rect 14850 80 14910 105
rect 14850 35 14905 80
rect 14905 35 14910 80
rect 15040 80 15100 105
rect 15040 35 15095 80
rect 15095 35 15100 80
rect 15235 80 15295 105
rect 15235 35 15290 80
rect 15290 35 15295 80
rect 15425 80 15485 105
rect 15425 35 15480 80
rect 15480 35 15485 80
rect 15620 80 15680 105
rect 15620 35 15675 80
rect 15675 35 15680 80
rect 15995 80 16055 105
rect 15995 35 16050 80
rect 16050 35 16055 80
rect 16185 80 16245 105
rect 16185 35 16240 80
rect 16240 35 16245 80
rect 16380 80 16440 105
rect 16380 35 16435 80
rect 16435 35 16440 80
rect 16575 80 16635 105
rect 16575 35 16630 80
rect 16630 35 16635 80
rect 16765 80 16825 105
rect 16765 35 16820 80
rect 16820 35 16825 80
rect 16960 80 17020 105
rect 16960 35 17015 80
rect 17015 35 17020 80
rect 17150 80 17210 105
rect 17150 35 17205 80
rect 17205 35 17210 80
rect 17345 80 17405 105
rect 17345 35 17400 80
rect 17400 35 17405 80
rect 17535 80 17595 105
rect 17535 35 17590 80
rect 17590 35 17595 80
rect 17725 80 17785 105
rect 17725 35 17780 80
rect 17780 35 17785 80
rect 17920 80 17980 105
rect 17920 35 17975 80
rect 17975 35 17980 80
rect 18110 80 18170 105
rect 18110 35 18165 80
rect 18165 35 18170 80
rect 18305 80 18365 105
rect 18305 35 18360 80
rect 18360 35 18365 80
rect 18495 80 18555 105
rect 18495 35 18550 80
rect 18550 35 18555 80
rect 18685 80 18745 105
rect 18685 35 18740 80
rect 18740 35 18745 80
rect 18880 80 18940 105
rect 18880 35 18935 80
rect 18935 35 18940 80
rect 19070 80 19130 105
rect 19070 35 19125 80
rect 19125 35 19130 80
rect 19265 80 19325 105
rect 19265 35 19320 80
rect 19320 35 19325 80
rect 19455 80 19515 105
rect 19455 35 19510 80
rect 19510 35 19515 80
rect 19645 80 19705 105
rect 19645 35 19700 80
rect 19700 35 19705 80
rect 19840 80 19900 105
rect 19840 35 19895 80
rect 19895 35 19900 80
rect 20030 80 20090 105
rect 20030 35 20085 80
rect 20085 35 20090 80
rect 20225 80 20285 105
rect 20225 35 20280 80
rect 20280 35 20285 80
rect 20415 80 20475 105
rect 20415 35 20470 80
rect 20470 35 20475 80
rect 20610 80 20670 105
rect 20610 35 20665 80
rect 20665 35 20670 80
rect 20800 80 20860 105
rect 20800 35 20855 80
rect 20855 35 20860 80
rect 20990 80 21050 105
rect 20990 35 21045 80
rect 21045 35 21050 80
rect 21185 80 21245 105
rect 21185 35 21240 80
rect 21240 35 21245 80
rect 21375 80 21435 105
rect 21375 35 21430 80
rect 21430 35 21435 80
rect 21565 80 21625 105
rect 21565 35 21620 80
rect 21620 35 21625 80
rect 21760 80 21820 105
rect 21760 35 21815 80
rect 21815 35 21820 80
rect 13795 -100 13850 -55
rect 13850 -100 13855 -55
rect 13795 -125 13855 -100
rect 13985 -100 14040 -55
rect 14040 -100 14045 -55
rect 13985 -125 14045 -100
rect 14180 -100 14235 -55
rect 14235 -100 14240 -55
rect 14180 -125 14240 -100
rect 14370 -100 14425 -55
rect 14425 -100 14430 -55
rect 14370 -125 14430 -100
rect 14560 -100 14615 -55
rect 14615 -100 14620 -55
rect 14560 -125 14620 -100
rect 14755 -100 14810 -55
rect 14810 -100 14815 -55
rect 14755 -125 14815 -100
rect 14945 -100 15000 -55
rect 15000 -100 15005 -55
rect 14945 -125 15005 -100
rect 15140 -100 15195 -55
rect 15195 -100 15200 -55
rect 15140 -125 15200 -100
rect 15330 -100 15385 -55
rect 15385 -100 15390 -55
rect 15330 -125 15390 -100
rect 15520 -100 15575 -55
rect 15575 -100 15580 -55
rect 15520 -125 15580 -100
rect 16090 -100 16095 -55
rect 16095 -100 16150 -55
rect 16090 -125 16150 -100
rect 16280 -100 16285 -55
rect 16285 -100 16340 -55
rect 16280 -125 16340 -100
rect 16475 -100 16480 -55
rect 16480 -100 16535 -55
rect 16475 -125 16535 -100
rect 16665 -100 16670 -55
rect 16670 -100 16725 -55
rect 16665 -125 16725 -100
rect 16860 -100 16865 -55
rect 16865 -100 16920 -55
rect 16860 -125 16920 -100
rect 17045 -100 17050 -55
rect 17050 -100 17105 -55
rect 17045 -125 17105 -100
rect 17245 -100 17250 -55
rect 17250 -100 17305 -55
rect 17245 -125 17305 -100
rect 17430 -100 17435 -55
rect 17435 -100 17490 -55
rect 17430 -125 17490 -100
rect 17625 -100 17630 -55
rect 17630 -100 17685 -55
rect 17625 -125 17685 -100
rect 17820 -100 17825 -55
rect 17825 -100 17880 -55
rect 17820 -125 17880 -100
rect 18005 -100 18010 -55
rect 18010 -100 18065 -55
rect 18005 -125 18065 -100
rect 18200 -100 18205 -55
rect 18205 -100 18260 -55
rect 18200 -125 18260 -100
rect 18390 -100 18395 -55
rect 18395 -100 18450 -55
rect 18390 -125 18450 -100
rect 18585 -100 18590 -55
rect 18590 -100 18645 -55
rect 18585 -125 18645 -100
rect 18775 -100 18780 -55
rect 18780 -100 18835 -55
rect 18775 -125 18835 -100
rect 18970 -100 18975 -55
rect 18975 -100 19030 -55
rect 18970 -125 19030 -100
rect 19160 -100 19165 -55
rect 19165 -100 19220 -55
rect 19160 -125 19220 -100
rect 19355 -100 19360 -55
rect 19360 -100 19415 -55
rect 19355 -125 19415 -100
rect 19545 -100 19550 -55
rect 19550 -100 19605 -55
rect 19545 -125 19605 -100
rect 19740 -100 19745 -55
rect 19745 -100 19800 -55
rect 19740 -125 19800 -100
rect 19930 -100 19935 -55
rect 19935 -100 19990 -55
rect 19930 -125 19990 -100
rect 20120 -100 20125 -55
rect 20125 -100 20180 -55
rect 20120 -125 20180 -100
rect 20315 -100 20320 -55
rect 20320 -100 20375 -55
rect 20315 -125 20375 -100
rect 20505 -100 20510 -55
rect 20510 -100 20565 -55
rect 20505 -125 20565 -100
rect 20700 -100 20705 -55
rect 20705 -100 20760 -55
rect 20700 -125 20760 -100
rect 20890 -100 20895 -55
rect 20895 -100 20950 -55
rect 20890 -125 20950 -100
rect 21080 -100 21085 -55
rect 21085 -100 21140 -55
rect 21080 -125 21140 -100
rect 21275 -100 21280 -55
rect 21280 -100 21335 -55
rect 21275 -125 21335 -100
rect 21465 -100 21470 -55
rect 21470 -100 21525 -55
rect 21465 -125 21525 -100
rect 21655 -100 21660 -55
rect 21660 -100 21715 -55
rect 21655 -125 21715 -100
rect 10205 -1080 10600 -550
rect 13750 -1655 14135 -560
rect 17460 -1655 17845 -565
<< metal3 >>
rect 13725 2320 14160 2475
rect 13715 2280 14160 2320
rect 10190 1720 10640 1735
rect 10190 1190 10210 1720
rect 10605 1190 10640 1720
rect 10190 -550 10640 1190
rect 13715 1190 13740 2280
rect 14120 2040 14160 2280
rect 17435 2280 17870 2310
rect 14120 1190 14150 2040
rect 13715 1090 14150 1190
rect 17435 1190 17455 2280
rect 17840 1190 17870 2280
rect 17435 1165 17870 1190
rect 13715 765 15710 1090
rect 13715 745 13795 765
rect 13785 695 13795 745
rect 13855 695 13985 765
rect 14045 695 14180 765
rect 14240 695 14370 765
rect 14430 695 14560 765
rect 14620 695 14755 765
rect 14815 695 14945 765
rect 15005 695 15140 765
rect 15200 695 15330 765
rect 15390 695 15520 765
rect 15580 695 15710 765
rect 13785 685 15710 695
rect 15980 765 22825 1100
rect 15980 695 16090 765
rect 16150 695 16280 765
rect 16340 695 16475 765
rect 16535 695 16665 765
rect 16725 695 16860 765
rect 16920 695 17045 765
rect 17105 695 17245 765
rect 17305 695 17430 765
rect 17490 695 17625 765
rect 17685 695 17820 765
rect 17880 695 18005 765
rect 18065 695 18200 765
rect 18260 695 18390 765
rect 18450 695 18585 765
rect 18645 695 18775 765
rect 18835 695 18970 765
rect 19030 695 19160 765
rect 19220 695 19355 765
rect 19415 695 19545 765
rect 19605 695 19740 765
rect 19800 695 19930 765
rect 19990 695 20120 765
rect 20180 695 20315 765
rect 20375 695 20505 765
rect 20565 695 20700 765
rect 20760 695 20890 765
rect 20950 695 21080 765
rect 21140 695 21275 765
rect 21335 695 21465 765
rect 21525 695 21655 765
rect 21715 695 21820 765
rect 15980 685 21820 695
rect 13680 605 21825 615
rect 13680 535 13700 605
rect 13760 535 13890 605
rect 13950 535 14085 605
rect 14145 535 14275 605
rect 14335 535 14470 605
rect 14530 535 14655 605
rect 14715 535 14850 605
rect 14910 535 15040 605
rect 15100 535 15235 605
rect 15295 535 15425 605
rect 15485 535 15620 605
rect 15680 535 15995 605
rect 16055 535 16185 605
rect 16245 535 16380 605
rect 16440 535 16575 605
rect 16635 535 16765 605
rect 16825 535 16960 605
rect 17020 535 17150 605
rect 17210 535 17345 605
rect 17405 535 17535 605
rect 17595 535 17725 605
rect 17785 535 17920 605
rect 17980 535 18110 605
rect 18170 535 18305 605
rect 18365 535 18495 605
rect 18555 535 18685 605
rect 18745 535 18880 605
rect 18940 535 19070 605
rect 19130 535 19265 605
rect 19325 535 19455 605
rect 19515 535 19645 605
rect 19705 535 19840 605
rect 19900 535 20030 605
rect 20090 535 20225 605
rect 20285 535 20415 605
rect 20475 535 20610 605
rect 20670 535 20800 605
rect 20860 535 20990 605
rect 21050 535 21185 605
rect 21245 535 21375 605
rect 21435 535 21565 605
rect 21625 535 21760 605
rect 21820 535 21825 605
rect 13680 105 21825 535
rect 13680 35 13700 105
rect 13760 35 13890 105
rect 13950 35 14085 105
rect 14145 35 14275 105
rect 14335 35 14470 105
rect 14530 35 14655 105
rect 14715 35 14850 105
rect 14910 35 15040 105
rect 15100 35 15235 105
rect 15295 35 15425 105
rect 15485 35 15620 105
rect 15680 35 15995 105
rect 16055 35 16185 105
rect 16245 35 16380 105
rect 16440 35 16575 105
rect 16635 35 16765 105
rect 16825 35 16960 105
rect 17020 35 17150 105
rect 17210 35 17345 105
rect 17405 35 17535 105
rect 17595 35 17725 105
rect 17785 35 17920 105
rect 17980 35 18110 105
rect 18170 35 18305 105
rect 18365 35 18495 105
rect 18555 35 18685 105
rect 18745 35 18880 105
rect 18940 35 19070 105
rect 19130 35 19265 105
rect 19325 35 19455 105
rect 19515 35 19645 105
rect 19705 35 19840 105
rect 19900 35 20030 105
rect 20090 35 20225 105
rect 20285 35 20415 105
rect 20475 35 20610 105
rect 20670 35 20800 105
rect 20860 35 20990 105
rect 21050 35 21185 105
rect 21245 35 21375 105
rect 21435 35 21565 105
rect 21625 35 21760 105
rect 21820 35 21825 105
rect 13680 25 21825 35
rect 22025 -45 22825 765
rect 10190 -1080 10205 -550
rect 10600 -1080 10640 -550
rect 10190 -1275 10640 -1080
rect 13725 -55 15710 -45
rect 13725 -125 13795 -55
rect 13855 -125 13985 -55
rect 14045 -125 14180 -55
rect 14240 -125 14370 -55
rect 14430 -125 14560 -55
rect 14620 -125 14755 -55
rect 14815 -125 14945 -55
rect 15005 -125 15140 -55
rect 15200 -125 15330 -55
rect 15390 -125 15520 -55
rect 15580 -125 15710 -55
rect 13725 -455 15710 -125
rect 15980 -55 22825 -45
rect 15980 -125 16090 -55
rect 16150 -125 16280 -55
rect 16340 -125 16475 -55
rect 16535 -125 16665 -55
rect 16725 -125 16860 -55
rect 16920 -125 17045 -55
rect 17105 -125 17245 -55
rect 17305 -125 17430 -55
rect 17490 -125 17625 -55
rect 17685 -125 17820 -55
rect 17880 -125 18005 -55
rect 18065 -125 18200 -55
rect 18260 -125 18390 -55
rect 18450 -125 18585 -55
rect 18645 -125 18775 -55
rect 18835 -125 18970 -55
rect 19030 -125 19160 -55
rect 19220 -125 19355 -55
rect 19415 -125 19545 -55
rect 19605 -125 19740 -55
rect 19800 -125 19930 -55
rect 19990 -125 20120 -55
rect 20180 -125 20315 -55
rect 20375 -125 20505 -55
rect 20565 -125 20700 -55
rect 20760 -125 20890 -55
rect 20950 -125 21080 -55
rect 21140 -125 21275 -55
rect 21335 -125 21465 -55
rect 21525 -125 21655 -55
rect 21715 -125 22825 -55
rect 15980 -455 22825 -125
rect 13725 -560 14160 -455
rect 13725 -1655 13750 -560
rect 14135 -1430 14160 -560
rect 17435 -565 17870 -530
rect 14135 -1655 14165 -1430
rect 13725 -1680 14165 -1655
rect 17435 -1655 17460 -565
rect 17845 -1655 17870 -565
rect 17435 -1675 17870 -1655
rect 13730 -1865 14165 -1680
rect 22025 -1795 22825 -455
<< via3 >>
rect 17455 1190 17840 2280
rect 17460 -1655 17845 -565
<< metal4 >>
rect 17435 2280 18025 2310
rect 17435 1190 17455 2280
rect 17840 1190 18025 2280
rect 17435 -565 18025 1190
rect 17435 -1655 17460 -565
rect 17845 -1655 18025 -565
rect 17435 -1675 18025 -1655
rect 17440 -1680 18025 -1675
use sky130_fd_pr__nfet_01v8_lvt_YTLFGX  XM1 
timestamp 1662510845
transform 1 0 10847 0 -1 650
box -1127 -310 1127 310
use sky130_fd_pr__nfet_01v8_lvt_YTLFGX  XM2
timestamp 1662510845
transform 1 0 10847 0 1 -10
box -1127 -310 1127 310
use sky130_fd_pr__nfet_01v8_lvt_LELFGX  XM3
timestamp 1662407989
transform 1 0 18902 0 1 650
box -3047 -310 3047 310
use sky130_fd_pr__nfet_01v8_lvt_LELFGX  XM4
timestamp 1662407989
transform 1 0 18902 0 1 -10
box -3047 -310 3047 310
use sky130_fd_pr__nfet_01v8_lvt_YTLFGX  XM32
timestamp 1662510845
transform 1 0 14687 0 1 650
box -1127 -310 1127 310
use sky130_fd_pr__nfet_01v8_lvt_YTLFGX  XM33
timestamp 1662510845
transform 1 0 14687 0 -1 -10
box -1127 -310 1127 310
use sky130_fd_pr__nfet_01v8_lvt_HNLS5R  XM42 
timestamp 1662515274
transform 1 0 12379 0 -1 650
box -359 -310 359 310
use sky130_fd_pr__nfet_01v8_lvt_HNLS5R  XM43
timestamp 1662515274
transform 1 0 12379 0 1 -10
box -359 -310 359 310
use sky130_fd_pr__res_high_po_2p85_P79JE3  XR1 
timestamp 1662404926
transform 0 1 11383 -1 0 1451
box -451 -1358 451 1358
use sky130_fd_pr__res_high_po_2p85_P79JE3  XR2
timestamp 1662404926
transform 0 1 11380 -1 0 -807
box -451 -1358 451 1358
use sky130_fd_pr__res_high_po_5p73_W59YBA  XR3
timestamp 1662407989
transform 0 1 15798 -1 0 -1101
box -739 -2238 739 2238
use sky130_fd_pr__res_high_po_5p73_W59YBA  XR29
timestamp 1662407989
transform 0 1 15798 -1 0 1739
box -739 -2238 739 2238
<< labels >>
rlabel metal1 11925 -1260 11975 830 1 BIAS
rlabel metal2 8845 -1300 9445 980 1 GND
rlabel metal3 10190 -1275 10640 -1080 1 VDD
rlabel metal1 12900 -1255 12955 175 1 INB
rlabel metal1 13365 -1260 13415 520 1 INA
rlabel metal3 22025 -1795 22825 -240 1 GND
rlabel metal4 17440 -1680 18025 2310 1 VDD
rlabel metal1 15855 -1840 15905 830 1 BIAS
rlabel locali 12675 1830 13610 1870 1 SUB
rlabel metal3 13725 2280 14160 2475 1 OUTA
rlabel metal3 13730 -1865 14165 -1655 1 OUTB
<< end >>
