magic
tech sky130A
magscale 1 2
timestamp 1662988209
<< error_p >>
rect -29 5815 29 5821
rect -29 5781 -17 5815
rect -29 5775 29 5781
rect -29 5505 29 5511
rect -29 5471 -17 5505
rect -29 5465 29 5471
rect -29 5397 29 5403
rect -29 5363 -17 5397
rect -29 5357 29 5363
rect -29 5087 29 5093
rect -29 5053 -17 5087
rect -29 5047 29 5053
rect -29 4979 29 4985
rect -29 4945 -17 4979
rect -29 4939 29 4945
rect -29 4669 29 4675
rect -29 4635 -17 4669
rect -29 4629 29 4635
rect -29 4561 29 4567
rect -29 4527 -17 4561
rect -29 4521 29 4527
rect -29 4251 29 4257
rect -29 4217 -17 4251
rect -29 4211 29 4217
rect -29 4143 29 4149
rect -29 4109 -17 4143
rect -29 4103 29 4109
rect -29 3833 29 3839
rect -29 3799 -17 3833
rect -29 3793 29 3799
rect -29 3725 29 3731
rect -29 3691 -17 3725
rect -29 3685 29 3691
rect -29 3415 29 3421
rect -29 3381 -17 3415
rect -29 3375 29 3381
rect -29 3307 29 3313
rect -29 3273 -17 3307
rect -29 3267 29 3273
rect -29 2997 29 3003
rect -29 2963 -17 2997
rect -29 2957 29 2963
rect -29 2889 29 2895
rect -29 2855 -17 2889
rect -29 2849 29 2855
rect -29 2579 29 2585
rect -29 2545 -17 2579
rect -29 2539 29 2545
rect -29 2471 29 2477
rect -29 2437 -17 2471
rect -29 2431 29 2437
rect -29 2161 29 2167
rect -29 2127 -17 2161
rect -29 2121 29 2127
rect -29 2053 29 2059
rect -29 2019 -17 2053
rect -29 2013 29 2019
rect -29 1743 29 1749
rect -29 1709 -17 1743
rect -29 1703 29 1709
rect -29 1635 29 1641
rect -29 1601 -17 1635
rect -29 1595 29 1601
rect -29 1325 29 1331
rect -29 1291 -17 1325
rect -29 1285 29 1291
rect -29 1217 29 1223
rect -29 1183 -17 1217
rect -29 1177 29 1183
rect -29 907 29 913
rect -29 873 -17 907
rect -29 867 29 873
rect -29 799 29 805
rect -29 765 -17 799
rect -29 759 29 765
rect -29 489 29 495
rect -29 455 -17 489
rect -29 449 29 455
rect -29 381 29 387
rect -29 347 -17 381
rect -29 341 29 347
rect -29 71 29 77
rect -29 37 -17 71
rect -29 31 29 37
rect -29 -37 29 -31
rect -29 -71 -17 -37
rect -29 -77 29 -71
rect -29 -347 29 -341
rect -29 -381 -17 -347
rect -29 -387 29 -381
rect -29 -455 29 -449
rect -29 -489 -17 -455
rect -29 -495 29 -489
rect -29 -765 29 -759
rect -29 -799 -17 -765
rect -29 -805 29 -799
rect -29 -873 29 -867
rect -29 -907 -17 -873
rect -29 -913 29 -907
rect -29 -1183 29 -1177
rect -29 -1217 -17 -1183
rect -29 -1223 29 -1217
rect -29 -1291 29 -1285
rect -29 -1325 -17 -1291
rect -29 -1331 29 -1325
rect -29 -1601 29 -1595
rect -29 -1635 -17 -1601
rect -29 -1641 29 -1635
rect -29 -1709 29 -1703
rect -29 -1743 -17 -1709
rect -29 -1749 29 -1743
rect -29 -2019 29 -2013
rect -29 -2053 -17 -2019
rect -29 -2059 29 -2053
rect -29 -2127 29 -2121
rect -29 -2161 -17 -2127
rect -29 -2167 29 -2161
rect -29 -2437 29 -2431
rect -29 -2471 -17 -2437
rect -29 -2477 29 -2471
rect -29 -2545 29 -2539
rect -29 -2579 -17 -2545
rect -29 -2585 29 -2579
rect -29 -2855 29 -2849
rect -29 -2889 -17 -2855
rect -29 -2895 29 -2889
rect -29 -2963 29 -2957
rect -29 -2997 -17 -2963
rect -29 -3003 29 -2997
rect -29 -3273 29 -3267
rect -29 -3307 -17 -3273
rect -29 -3313 29 -3307
rect -29 -3381 29 -3375
rect -29 -3415 -17 -3381
rect -29 -3421 29 -3415
rect -29 -3691 29 -3685
rect -29 -3725 -17 -3691
rect -29 -3731 29 -3725
rect -29 -3799 29 -3793
rect -29 -3833 -17 -3799
rect -29 -3839 29 -3833
rect -29 -4109 29 -4103
rect -29 -4143 -17 -4109
rect -29 -4149 29 -4143
rect -29 -4217 29 -4211
rect -29 -4251 -17 -4217
rect -29 -4257 29 -4251
rect -29 -4527 29 -4521
rect -29 -4561 -17 -4527
rect -29 -4567 29 -4561
rect -29 -4635 29 -4629
rect -29 -4669 -17 -4635
rect -29 -4675 29 -4669
rect -29 -4945 29 -4939
rect -29 -4979 -17 -4945
rect -29 -4985 29 -4979
rect -29 -5053 29 -5047
rect -29 -5087 -17 -5053
rect -29 -5093 29 -5087
rect -29 -5363 29 -5357
rect -29 -5397 -17 -5363
rect -29 -5403 29 -5397
rect -29 -5471 29 -5465
rect -29 -5505 -17 -5471
rect -29 -5511 29 -5505
rect -29 -5781 29 -5775
rect -29 -5815 -17 -5781
rect -29 -5821 29 -5815
<< pwell >>
rect -211 -5953 211 5953
<< nmoslvt >>
rect -15 5543 15 5743
rect -15 5125 15 5325
rect -15 4707 15 4907
rect -15 4289 15 4489
rect -15 3871 15 4071
rect -15 3453 15 3653
rect -15 3035 15 3235
rect -15 2617 15 2817
rect -15 2199 15 2399
rect -15 1781 15 1981
rect -15 1363 15 1563
rect -15 945 15 1145
rect -15 527 15 727
rect -15 109 15 309
rect -15 -309 15 -109
rect -15 -727 15 -527
rect -15 -1145 15 -945
rect -15 -1563 15 -1363
rect -15 -1981 15 -1781
rect -15 -2399 15 -2199
rect -15 -2817 15 -2617
rect -15 -3235 15 -3035
rect -15 -3653 15 -3453
rect -15 -4071 15 -3871
rect -15 -4489 15 -4289
rect -15 -4907 15 -4707
rect -15 -5325 15 -5125
rect -15 -5743 15 -5543
<< ndiff >>
rect -73 5731 -15 5743
rect -73 5555 -61 5731
rect -27 5555 -15 5731
rect -73 5543 -15 5555
rect 15 5731 73 5743
rect 15 5555 27 5731
rect 61 5555 73 5731
rect 15 5543 73 5555
rect -73 5313 -15 5325
rect -73 5137 -61 5313
rect -27 5137 -15 5313
rect -73 5125 -15 5137
rect 15 5313 73 5325
rect 15 5137 27 5313
rect 61 5137 73 5313
rect 15 5125 73 5137
rect -73 4895 -15 4907
rect -73 4719 -61 4895
rect -27 4719 -15 4895
rect -73 4707 -15 4719
rect 15 4895 73 4907
rect 15 4719 27 4895
rect 61 4719 73 4895
rect 15 4707 73 4719
rect -73 4477 -15 4489
rect -73 4301 -61 4477
rect -27 4301 -15 4477
rect -73 4289 -15 4301
rect 15 4477 73 4489
rect 15 4301 27 4477
rect 61 4301 73 4477
rect 15 4289 73 4301
rect -73 4059 -15 4071
rect -73 3883 -61 4059
rect -27 3883 -15 4059
rect -73 3871 -15 3883
rect 15 4059 73 4071
rect 15 3883 27 4059
rect 61 3883 73 4059
rect 15 3871 73 3883
rect -73 3641 -15 3653
rect -73 3465 -61 3641
rect -27 3465 -15 3641
rect -73 3453 -15 3465
rect 15 3641 73 3653
rect 15 3465 27 3641
rect 61 3465 73 3641
rect 15 3453 73 3465
rect -73 3223 -15 3235
rect -73 3047 -61 3223
rect -27 3047 -15 3223
rect -73 3035 -15 3047
rect 15 3223 73 3235
rect 15 3047 27 3223
rect 61 3047 73 3223
rect 15 3035 73 3047
rect -73 2805 -15 2817
rect -73 2629 -61 2805
rect -27 2629 -15 2805
rect -73 2617 -15 2629
rect 15 2805 73 2817
rect 15 2629 27 2805
rect 61 2629 73 2805
rect 15 2617 73 2629
rect -73 2387 -15 2399
rect -73 2211 -61 2387
rect -27 2211 -15 2387
rect -73 2199 -15 2211
rect 15 2387 73 2399
rect 15 2211 27 2387
rect 61 2211 73 2387
rect 15 2199 73 2211
rect -73 1969 -15 1981
rect -73 1793 -61 1969
rect -27 1793 -15 1969
rect -73 1781 -15 1793
rect 15 1969 73 1981
rect 15 1793 27 1969
rect 61 1793 73 1969
rect 15 1781 73 1793
rect -73 1551 -15 1563
rect -73 1375 -61 1551
rect -27 1375 -15 1551
rect -73 1363 -15 1375
rect 15 1551 73 1563
rect 15 1375 27 1551
rect 61 1375 73 1551
rect 15 1363 73 1375
rect -73 1133 -15 1145
rect -73 957 -61 1133
rect -27 957 -15 1133
rect -73 945 -15 957
rect 15 1133 73 1145
rect 15 957 27 1133
rect 61 957 73 1133
rect 15 945 73 957
rect -73 715 -15 727
rect -73 539 -61 715
rect -27 539 -15 715
rect -73 527 -15 539
rect 15 715 73 727
rect 15 539 27 715
rect 61 539 73 715
rect 15 527 73 539
rect -73 297 -15 309
rect -73 121 -61 297
rect -27 121 -15 297
rect -73 109 -15 121
rect 15 297 73 309
rect 15 121 27 297
rect 61 121 73 297
rect 15 109 73 121
rect -73 -121 -15 -109
rect -73 -297 -61 -121
rect -27 -297 -15 -121
rect -73 -309 -15 -297
rect 15 -121 73 -109
rect 15 -297 27 -121
rect 61 -297 73 -121
rect 15 -309 73 -297
rect -73 -539 -15 -527
rect -73 -715 -61 -539
rect -27 -715 -15 -539
rect -73 -727 -15 -715
rect 15 -539 73 -527
rect 15 -715 27 -539
rect 61 -715 73 -539
rect 15 -727 73 -715
rect -73 -957 -15 -945
rect -73 -1133 -61 -957
rect -27 -1133 -15 -957
rect -73 -1145 -15 -1133
rect 15 -957 73 -945
rect 15 -1133 27 -957
rect 61 -1133 73 -957
rect 15 -1145 73 -1133
rect -73 -1375 -15 -1363
rect -73 -1551 -61 -1375
rect -27 -1551 -15 -1375
rect -73 -1563 -15 -1551
rect 15 -1375 73 -1363
rect 15 -1551 27 -1375
rect 61 -1551 73 -1375
rect 15 -1563 73 -1551
rect -73 -1793 -15 -1781
rect -73 -1969 -61 -1793
rect -27 -1969 -15 -1793
rect -73 -1981 -15 -1969
rect 15 -1793 73 -1781
rect 15 -1969 27 -1793
rect 61 -1969 73 -1793
rect 15 -1981 73 -1969
rect -73 -2211 -15 -2199
rect -73 -2387 -61 -2211
rect -27 -2387 -15 -2211
rect -73 -2399 -15 -2387
rect 15 -2211 73 -2199
rect 15 -2387 27 -2211
rect 61 -2387 73 -2211
rect 15 -2399 73 -2387
rect -73 -2629 -15 -2617
rect -73 -2805 -61 -2629
rect -27 -2805 -15 -2629
rect -73 -2817 -15 -2805
rect 15 -2629 73 -2617
rect 15 -2805 27 -2629
rect 61 -2805 73 -2629
rect 15 -2817 73 -2805
rect -73 -3047 -15 -3035
rect -73 -3223 -61 -3047
rect -27 -3223 -15 -3047
rect -73 -3235 -15 -3223
rect 15 -3047 73 -3035
rect 15 -3223 27 -3047
rect 61 -3223 73 -3047
rect 15 -3235 73 -3223
rect -73 -3465 -15 -3453
rect -73 -3641 -61 -3465
rect -27 -3641 -15 -3465
rect -73 -3653 -15 -3641
rect 15 -3465 73 -3453
rect 15 -3641 27 -3465
rect 61 -3641 73 -3465
rect 15 -3653 73 -3641
rect -73 -3883 -15 -3871
rect -73 -4059 -61 -3883
rect -27 -4059 -15 -3883
rect -73 -4071 -15 -4059
rect 15 -3883 73 -3871
rect 15 -4059 27 -3883
rect 61 -4059 73 -3883
rect 15 -4071 73 -4059
rect -73 -4301 -15 -4289
rect -73 -4477 -61 -4301
rect -27 -4477 -15 -4301
rect -73 -4489 -15 -4477
rect 15 -4301 73 -4289
rect 15 -4477 27 -4301
rect 61 -4477 73 -4301
rect 15 -4489 73 -4477
rect -73 -4719 -15 -4707
rect -73 -4895 -61 -4719
rect -27 -4895 -15 -4719
rect -73 -4907 -15 -4895
rect 15 -4719 73 -4707
rect 15 -4895 27 -4719
rect 61 -4895 73 -4719
rect 15 -4907 73 -4895
rect -73 -5137 -15 -5125
rect -73 -5313 -61 -5137
rect -27 -5313 -15 -5137
rect -73 -5325 -15 -5313
rect 15 -5137 73 -5125
rect 15 -5313 27 -5137
rect 61 -5313 73 -5137
rect 15 -5325 73 -5313
rect -73 -5555 -15 -5543
rect -73 -5731 -61 -5555
rect -27 -5731 -15 -5555
rect -73 -5743 -15 -5731
rect 15 -5555 73 -5543
rect 15 -5731 27 -5555
rect 61 -5731 73 -5555
rect 15 -5743 73 -5731
<< ndiffc >>
rect -61 5555 -27 5731
rect 27 5555 61 5731
rect -61 5137 -27 5313
rect 27 5137 61 5313
rect -61 4719 -27 4895
rect 27 4719 61 4895
rect -61 4301 -27 4477
rect 27 4301 61 4477
rect -61 3883 -27 4059
rect 27 3883 61 4059
rect -61 3465 -27 3641
rect 27 3465 61 3641
rect -61 3047 -27 3223
rect 27 3047 61 3223
rect -61 2629 -27 2805
rect 27 2629 61 2805
rect -61 2211 -27 2387
rect 27 2211 61 2387
rect -61 1793 -27 1969
rect 27 1793 61 1969
rect -61 1375 -27 1551
rect 27 1375 61 1551
rect -61 957 -27 1133
rect 27 957 61 1133
rect -61 539 -27 715
rect 27 539 61 715
rect -61 121 -27 297
rect 27 121 61 297
rect -61 -297 -27 -121
rect 27 -297 61 -121
rect -61 -715 -27 -539
rect 27 -715 61 -539
rect -61 -1133 -27 -957
rect 27 -1133 61 -957
rect -61 -1551 -27 -1375
rect 27 -1551 61 -1375
rect -61 -1969 -27 -1793
rect 27 -1969 61 -1793
rect -61 -2387 -27 -2211
rect 27 -2387 61 -2211
rect -61 -2805 -27 -2629
rect 27 -2805 61 -2629
rect -61 -3223 -27 -3047
rect 27 -3223 61 -3047
rect -61 -3641 -27 -3465
rect 27 -3641 61 -3465
rect -61 -4059 -27 -3883
rect 27 -4059 61 -3883
rect -61 -4477 -27 -4301
rect 27 -4477 61 -4301
rect -61 -4895 -27 -4719
rect 27 -4895 61 -4719
rect -61 -5313 -27 -5137
rect 27 -5313 61 -5137
rect -61 -5731 -27 -5555
rect 27 -5731 61 -5555
<< psubdiff >>
rect -175 5883 -79 5917
rect 79 5883 175 5917
rect -175 5821 -141 5883
rect 141 5821 175 5883
rect -175 -5883 -141 -5821
rect 141 -5883 175 -5821
rect -175 -5917 -79 -5883
rect 79 -5917 175 -5883
<< psubdiffcont >>
rect -79 5883 79 5917
rect -175 -5821 -141 5821
rect 141 -5821 175 5821
rect -79 -5917 79 -5883
<< poly >>
rect -33 5815 33 5831
rect -33 5781 -17 5815
rect 17 5781 33 5815
rect -33 5765 33 5781
rect -15 5743 15 5765
rect -15 5521 15 5543
rect -33 5505 33 5521
rect -33 5471 -17 5505
rect 17 5471 33 5505
rect -33 5455 33 5471
rect -33 5397 33 5413
rect -33 5363 -17 5397
rect 17 5363 33 5397
rect -33 5347 33 5363
rect -15 5325 15 5347
rect -15 5103 15 5125
rect -33 5087 33 5103
rect -33 5053 -17 5087
rect 17 5053 33 5087
rect -33 5037 33 5053
rect -33 4979 33 4995
rect -33 4945 -17 4979
rect 17 4945 33 4979
rect -33 4929 33 4945
rect -15 4907 15 4929
rect -15 4685 15 4707
rect -33 4669 33 4685
rect -33 4635 -17 4669
rect 17 4635 33 4669
rect -33 4619 33 4635
rect -33 4561 33 4577
rect -33 4527 -17 4561
rect 17 4527 33 4561
rect -33 4511 33 4527
rect -15 4489 15 4511
rect -15 4267 15 4289
rect -33 4251 33 4267
rect -33 4217 -17 4251
rect 17 4217 33 4251
rect -33 4201 33 4217
rect -33 4143 33 4159
rect -33 4109 -17 4143
rect 17 4109 33 4143
rect -33 4093 33 4109
rect -15 4071 15 4093
rect -15 3849 15 3871
rect -33 3833 33 3849
rect -33 3799 -17 3833
rect 17 3799 33 3833
rect -33 3783 33 3799
rect -33 3725 33 3741
rect -33 3691 -17 3725
rect 17 3691 33 3725
rect -33 3675 33 3691
rect -15 3653 15 3675
rect -15 3431 15 3453
rect -33 3415 33 3431
rect -33 3381 -17 3415
rect 17 3381 33 3415
rect -33 3365 33 3381
rect -33 3307 33 3323
rect -33 3273 -17 3307
rect 17 3273 33 3307
rect -33 3257 33 3273
rect -15 3235 15 3257
rect -15 3013 15 3035
rect -33 2997 33 3013
rect -33 2963 -17 2997
rect 17 2963 33 2997
rect -33 2947 33 2963
rect -33 2889 33 2905
rect -33 2855 -17 2889
rect 17 2855 33 2889
rect -33 2839 33 2855
rect -15 2817 15 2839
rect -15 2595 15 2617
rect -33 2579 33 2595
rect -33 2545 -17 2579
rect 17 2545 33 2579
rect -33 2529 33 2545
rect -33 2471 33 2487
rect -33 2437 -17 2471
rect 17 2437 33 2471
rect -33 2421 33 2437
rect -15 2399 15 2421
rect -15 2177 15 2199
rect -33 2161 33 2177
rect -33 2127 -17 2161
rect 17 2127 33 2161
rect -33 2111 33 2127
rect -33 2053 33 2069
rect -33 2019 -17 2053
rect 17 2019 33 2053
rect -33 2003 33 2019
rect -15 1981 15 2003
rect -15 1759 15 1781
rect -33 1743 33 1759
rect -33 1709 -17 1743
rect 17 1709 33 1743
rect -33 1693 33 1709
rect -33 1635 33 1651
rect -33 1601 -17 1635
rect 17 1601 33 1635
rect -33 1585 33 1601
rect -15 1563 15 1585
rect -15 1341 15 1363
rect -33 1325 33 1341
rect -33 1291 -17 1325
rect 17 1291 33 1325
rect -33 1275 33 1291
rect -33 1217 33 1233
rect -33 1183 -17 1217
rect 17 1183 33 1217
rect -33 1167 33 1183
rect -15 1145 15 1167
rect -15 923 15 945
rect -33 907 33 923
rect -33 873 -17 907
rect 17 873 33 907
rect -33 857 33 873
rect -33 799 33 815
rect -33 765 -17 799
rect 17 765 33 799
rect -33 749 33 765
rect -15 727 15 749
rect -15 505 15 527
rect -33 489 33 505
rect -33 455 -17 489
rect 17 455 33 489
rect -33 439 33 455
rect -33 381 33 397
rect -33 347 -17 381
rect 17 347 33 381
rect -33 331 33 347
rect -15 309 15 331
rect -15 87 15 109
rect -33 71 33 87
rect -33 37 -17 71
rect 17 37 33 71
rect -33 21 33 37
rect -33 -37 33 -21
rect -33 -71 -17 -37
rect 17 -71 33 -37
rect -33 -87 33 -71
rect -15 -109 15 -87
rect -15 -331 15 -309
rect -33 -347 33 -331
rect -33 -381 -17 -347
rect 17 -381 33 -347
rect -33 -397 33 -381
rect -33 -455 33 -439
rect -33 -489 -17 -455
rect 17 -489 33 -455
rect -33 -505 33 -489
rect -15 -527 15 -505
rect -15 -749 15 -727
rect -33 -765 33 -749
rect -33 -799 -17 -765
rect 17 -799 33 -765
rect -33 -815 33 -799
rect -33 -873 33 -857
rect -33 -907 -17 -873
rect 17 -907 33 -873
rect -33 -923 33 -907
rect -15 -945 15 -923
rect -15 -1167 15 -1145
rect -33 -1183 33 -1167
rect -33 -1217 -17 -1183
rect 17 -1217 33 -1183
rect -33 -1233 33 -1217
rect -33 -1291 33 -1275
rect -33 -1325 -17 -1291
rect 17 -1325 33 -1291
rect -33 -1341 33 -1325
rect -15 -1363 15 -1341
rect -15 -1585 15 -1563
rect -33 -1601 33 -1585
rect -33 -1635 -17 -1601
rect 17 -1635 33 -1601
rect -33 -1651 33 -1635
rect -33 -1709 33 -1693
rect -33 -1743 -17 -1709
rect 17 -1743 33 -1709
rect -33 -1759 33 -1743
rect -15 -1781 15 -1759
rect -15 -2003 15 -1981
rect -33 -2019 33 -2003
rect -33 -2053 -17 -2019
rect 17 -2053 33 -2019
rect -33 -2069 33 -2053
rect -33 -2127 33 -2111
rect -33 -2161 -17 -2127
rect 17 -2161 33 -2127
rect -33 -2177 33 -2161
rect -15 -2199 15 -2177
rect -15 -2421 15 -2399
rect -33 -2437 33 -2421
rect -33 -2471 -17 -2437
rect 17 -2471 33 -2437
rect -33 -2487 33 -2471
rect -33 -2545 33 -2529
rect -33 -2579 -17 -2545
rect 17 -2579 33 -2545
rect -33 -2595 33 -2579
rect -15 -2617 15 -2595
rect -15 -2839 15 -2817
rect -33 -2855 33 -2839
rect -33 -2889 -17 -2855
rect 17 -2889 33 -2855
rect -33 -2905 33 -2889
rect -33 -2963 33 -2947
rect -33 -2997 -17 -2963
rect 17 -2997 33 -2963
rect -33 -3013 33 -2997
rect -15 -3035 15 -3013
rect -15 -3257 15 -3235
rect -33 -3273 33 -3257
rect -33 -3307 -17 -3273
rect 17 -3307 33 -3273
rect -33 -3323 33 -3307
rect -33 -3381 33 -3365
rect -33 -3415 -17 -3381
rect 17 -3415 33 -3381
rect -33 -3431 33 -3415
rect -15 -3453 15 -3431
rect -15 -3675 15 -3653
rect -33 -3691 33 -3675
rect -33 -3725 -17 -3691
rect 17 -3725 33 -3691
rect -33 -3741 33 -3725
rect -33 -3799 33 -3783
rect -33 -3833 -17 -3799
rect 17 -3833 33 -3799
rect -33 -3849 33 -3833
rect -15 -3871 15 -3849
rect -15 -4093 15 -4071
rect -33 -4109 33 -4093
rect -33 -4143 -17 -4109
rect 17 -4143 33 -4109
rect -33 -4159 33 -4143
rect -33 -4217 33 -4201
rect -33 -4251 -17 -4217
rect 17 -4251 33 -4217
rect -33 -4267 33 -4251
rect -15 -4289 15 -4267
rect -15 -4511 15 -4489
rect -33 -4527 33 -4511
rect -33 -4561 -17 -4527
rect 17 -4561 33 -4527
rect -33 -4577 33 -4561
rect -33 -4635 33 -4619
rect -33 -4669 -17 -4635
rect 17 -4669 33 -4635
rect -33 -4685 33 -4669
rect -15 -4707 15 -4685
rect -15 -4929 15 -4907
rect -33 -4945 33 -4929
rect -33 -4979 -17 -4945
rect 17 -4979 33 -4945
rect -33 -4995 33 -4979
rect -33 -5053 33 -5037
rect -33 -5087 -17 -5053
rect 17 -5087 33 -5053
rect -33 -5103 33 -5087
rect -15 -5125 15 -5103
rect -15 -5347 15 -5325
rect -33 -5363 33 -5347
rect -33 -5397 -17 -5363
rect 17 -5397 33 -5363
rect -33 -5413 33 -5397
rect -33 -5471 33 -5455
rect -33 -5505 -17 -5471
rect 17 -5505 33 -5471
rect -33 -5521 33 -5505
rect -15 -5543 15 -5521
rect -15 -5765 15 -5743
rect -33 -5781 33 -5765
rect -33 -5815 -17 -5781
rect 17 -5815 33 -5781
rect -33 -5831 33 -5815
<< polycont >>
rect -17 5781 17 5815
rect -17 5471 17 5505
rect -17 5363 17 5397
rect -17 5053 17 5087
rect -17 4945 17 4979
rect -17 4635 17 4669
rect -17 4527 17 4561
rect -17 4217 17 4251
rect -17 4109 17 4143
rect -17 3799 17 3833
rect -17 3691 17 3725
rect -17 3381 17 3415
rect -17 3273 17 3307
rect -17 2963 17 2997
rect -17 2855 17 2889
rect -17 2545 17 2579
rect -17 2437 17 2471
rect -17 2127 17 2161
rect -17 2019 17 2053
rect -17 1709 17 1743
rect -17 1601 17 1635
rect -17 1291 17 1325
rect -17 1183 17 1217
rect -17 873 17 907
rect -17 765 17 799
rect -17 455 17 489
rect -17 347 17 381
rect -17 37 17 71
rect -17 -71 17 -37
rect -17 -381 17 -347
rect -17 -489 17 -455
rect -17 -799 17 -765
rect -17 -907 17 -873
rect -17 -1217 17 -1183
rect -17 -1325 17 -1291
rect -17 -1635 17 -1601
rect -17 -1743 17 -1709
rect -17 -2053 17 -2019
rect -17 -2161 17 -2127
rect -17 -2471 17 -2437
rect -17 -2579 17 -2545
rect -17 -2889 17 -2855
rect -17 -2997 17 -2963
rect -17 -3307 17 -3273
rect -17 -3415 17 -3381
rect -17 -3725 17 -3691
rect -17 -3833 17 -3799
rect -17 -4143 17 -4109
rect -17 -4251 17 -4217
rect -17 -4561 17 -4527
rect -17 -4669 17 -4635
rect -17 -4979 17 -4945
rect -17 -5087 17 -5053
rect -17 -5397 17 -5363
rect -17 -5505 17 -5471
rect -17 -5815 17 -5781
<< locali >>
rect -175 5883 -79 5917
rect 79 5883 175 5917
rect -175 5821 -141 5883
rect 141 5821 175 5883
rect -33 5781 -17 5815
rect 17 5781 33 5815
rect -61 5731 -27 5747
rect -61 5539 -27 5555
rect 27 5731 61 5747
rect 27 5539 61 5555
rect -33 5471 -17 5505
rect 17 5471 33 5505
rect -33 5363 -17 5397
rect 17 5363 33 5397
rect -61 5313 -27 5329
rect -61 5121 -27 5137
rect 27 5313 61 5329
rect 27 5121 61 5137
rect -33 5053 -17 5087
rect 17 5053 33 5087
rect -33 4945 -17 4979
rect 17 4945 33 4979
rect -61 4895 -27 4911
rect -61 4703 -27 4719
rect 27 4895 61 4911
rect 27 4703 61 4719
rect -33 4635 -17 4669
rect 17 4635 33 4669
rect -33 4527 -17 4561
rect 17 4527 33 4561
rect -61 4477 -27 4493
rect -61 4285 -27 4301
rect 27 4477 61 4493
rect 27 4285 61 4301
rect -33 4217 -17 4251
rect 17 4217 33 4251
rect -33 4109 -17 4143
rect 17 4109 33 4143
rect -61 4059 -27 4075
rect -61 3867 -27 3883
rect 27 4059 61 4075
rect 27 3867 61 3883
rect -33 3799 -17 3833
rect 17 3799 33 3833
rect -33 3691 -17 3725
rect 17 3691 33 3725
rect -61 3641 -27 3657
rect -61 3449 -27 3465
rect 27 3641 61 3657
rect 27 3449 61 3465
rect -33 3381 -17 3415
rect 17 3381 33 3415
rect -33 3273 -17 3307
rect 17 3273 33 3307
rect -61 3223 -27 3239
rect -61 3031 -27 3047
rect 27 3223 61 3239
rect 27 3031 61 3047
rect -33 2963 -17 2997
rect 17 2963 33 2997
rect -33 2855 -17 2889
rect 17 2855 33 2889
rect -61 2805 -27 2821
rect -61 2613 -27 2629
rect 27 2805 61 2821
rect 27 2613 61 2629
rect -33 2545 -17 2579
rect 17 2545 33 2579
rect -33 2437 -17 2471
rect 17 2437 33 2471
rect -61 2387 -27 2403
rect -61 2195 -27 2211
rect 27 2387 61 2403
rect 27 2195 61 2211
rect -33 2127 -17 2161
rect 17 2127 33 2161
rect -33 2019 -17 2053
rect 17 2019 33 2053
rect -61 1969 -27 1985
rect -61 1777 -27 1793
rect 27 1969 61 1985
rect 27 1777 61 1793
rect -33 1709 -17 1743
rect 17 1709 33 1743
rect -33 1601 -17 1635
rect 17 1601 33 1635
rect -61 1551 -27 1567
rect -61 1359 -27 1375
rect 27 1551 61 1567
rect 27 1359 61 1375
rect -33 1291 -17 1325
rect 17 1291 33 1325
rect -33 1183 -17 1217
rect 17 1183 33 1217
rect -61 1133 -27 1149
rect -61 941 -27 957
rect 27 1133 61 1149
rect 27 941 61 957
rect -33 873 -17 907
rect 17 873 33 907
rect -33 765 -17 799
rect 17 765 33 799
rect -61 715 -27 731
rect -61 523 -27 539
rect 27 715 61 731
rect 27 523 61 539
rect -33 455 -17 489
rect 17 455 33 489
rect -33 347 -17 381
rect 17 347 33 381
rect -61 297 -27 313
rect -61 105 -27 121
rect 27 297 61 313
rect 27 105 61 121
rect -33 37 -17 71
rect 17 37 33 71
rect -33 -71 -17 -37
rect 17 -71 33 -37
rect -61 -121 -27 -105
rect -61 -313 -27 -297
rect 27 -121 61 -105
rect 27 -313 61 -297
rect -33 -381 -17 -347
rect 17 -381 33 -347
rect -33 -489 -17 -455
rect 17 -489 33 -455
rect -61 -539 -27 -523
rect -61 -731 -27 -715
rect 27 -539 61 -523
rect 27 -731 61 -715
rect -33 -799 -17 -765
rect 17 -799 33 -765
rect -33 -907 -17 -873
rect 17 -907 33 -873
rect -61 -957 -27 -941
rect -61 -1149 -27 -1133
rect 27 -957 61 -941
rect 27 -1149 61 -1133
rect -33 -1217 -17 -1183
rect 17 -1217 33 -1183
rect -33 -1325 -17 -1291
rect 17 -1325 33 -1291
rect -61 -1375 -27 -1359
rect -61 -1567 -27 -1551
rect 27 -1375 61 -1359
rect 27 -1567 61 -1551
rect -33 -1635 -17 -1601
rect 17 -1635 33 -1601
rect -33 -1743 -17 -1709
rect 17 -1743 33 -1709
rect -61 -1793 -27 -1777
rect -61 -1985 -27 -1969
rect 27 -1793 61 -1777
rect 27 -1985 61 -1969
rect -33 -2053 -17 -2019
rect 17 -2053 33 -2019
rect -33 -2161 -17 -2127
rect 17 -2161 33 -2127
rect -61 -2211 -27 -2195
rect -61 -2403 -27 -2387
rect 27 -2211 61 -2195
rect 27 -2403 61 -2387
rect -33 -2471 -17 -2437
rect 17 -2471 33 -2437
rect -33 -2579 -17 -2545
rect 17 -2579 33 -2545
rect -61 -2629 -27 -2613
rect -61 -2821 -27 -2805
rect 27 -2629 61 -2613
rect 27 -2821 61 -2805
rect -33 -2889 -17 -2855
rect 17 -2889 33 -2855
rect -33 -2997 -17 -2963
rect 17 -2997 33 -2963
rect -61 -3047 -27 -3031
rect -61 -3239 -27 -3223
rect 27 -3047 61 -3031
rect 27 -3239 61 -3223
rect -33 -3307 -17 -3273
rect 17 -3307 33 -3273
rect -33 -3415 -17 -3381
rect 17 -3415 33 -3381
rect -61 -3465 -27 -3449
rect -61 -3657 -27 -3641
rect 27 -3465 61 -3449
rect 27 -3657 61 -3641
rect -33 -3725 -17 -3691
rect 17 -3725 33 -3691
rect -33 -3833 -17 -3799
rect 17 -3833 33 -3799
rect -61 -3883 -27 -3867
rect -61 -4075 -27 -4059
rect 27 -3883 61 -3867
rect 27 -4075 61 -4059
rect -33 -4143 -17 -4109
rect 17 -4143 33 -4109
rect -33 -4251 -17 -4217
rect 17 -4251 33 -4217
rect -61 -4301 -27 -4285
rect -61 -4493 -27 -4477
rect 27 -4301 61 -4285
rect 27 -4493 61 -4477
rect -33 -4561 -17 -4527
rect 17 -4561 33 -4527
rect -33 -4669 -17 -4635
rect 17 -4669 33 -4635
rect -61 -4719 -27 -4703
rect -61 -4911 -27 -4895
rect 27 -4719 61 -4703
rect 27 -4911 61 -4895
rect -33 -4979 -17 -4945
rect 17 -4979 33 -4945
rect -33 -5087 -17 -5053
rect 17 -5087 33 -5053
rect -61 -5137 -27 -5121
rect -61 -5329 -27 -5313
rect 27 -5137 61 -5121
rect 27 -5329 61 -5313
rect -33 -5397 -17 -5363
rect 17 -5397 33 -5363
rect -33 -5505 -17 -5471
rect 17 -5505 33 -5471
rect -61 -5555 -27 -5539
rect -61 -5747 -27 -5731
rect 27 -5555 61 -5539
rect 27 -5747 61 -5731
rect -33 -5815 -17 -5781
rect 17 -5815 33 -5781
rect -175 -5883 -141 -5821
rect 141 -5883 175 -5821
rect -175 -5917 -79 -5883
rect 79 -5917 175 -5883
<< viali >>
rect -17 5781 17 5815
rect -61 5555 -27 5731
rect 27 5555 61 5731
rect -17 5471 17 5505
rect -17 5363 17 5397
rect -61 5137 -27 5313
rect 27 5137 61 5313
rect -17 5053 17 5087
rect -17 4945 17 4979
rect -61 4719 -27 4895
rect 27 4719 61 4895
rect -17 4635 17 4669
rect -17 4527 17 4561
rect -61 4301 -27 4477
rect 27 4301 61 4477
rect -17 4217 17 4251
rect -17 4109 17 4143
rect -61 3883 -27 4059
rect 27 3883 61 4059
rect -17 3799 17 3833
rect -17 3691 17 3725
rect -61 3465 -27 3641
rect 27 3465 61 3641
rect -17 3381 17 3415
rect -17 3273 17 3307
rect -61 3047 -27 3223
rect 27 3047 61 3223
rect -17 2963 17 2997
rect -17 2855 17 2889
rect -61 2629 -27 2805
rect 27 2629 61 2805
rect -17 2545 17 2579
rect -17 2437 17 2471
rect -61 2211 -27 2387
rect 27 2211 61 2387
rect -17 2127 17 2161
rect -17 2019 17 2053
rect -61 1793 -27 1969
rect 27 1793 61 1969
rect -17 1709 17 1743
rect -17 1601 17 1635
rect -61 1375 -27 1551
rect 27 1375 61 1551
rect -17 1291 17 1325
rect -17 1183 17 1217
rect -61 957 -27 1133
rect 27 957 61 1133
rect -17 873 17 907
rect -17 765 17 799
rect -61 539 -27 715
rect 27 539 61 715
rect -17 455 17 489
rect -17 347 17 381
rect -61 121 -27 297
rect 27 121 61 297
rect -17 37 17 71
rect -17 -71 17 -37
rect -61 -297 -27 -121
rect 27 -297 61 -121
rect -17 -381 17 -347
rect -17 -489 17 -455
rect -61 -715 -27 -539
rect 27 -715 61 -539
rect -17 -799 17 -765
rect -17 -907 17 -873
rect -61 -1133 -27 -957
rect 27 -1133 61 -957
rect -17 -1217 17 -1183
rect -17 -1325 17 -1291
rect -61 -1551 -27 -1375
rect 27 -1551 61 -1375
rect -17 -1635 17 -1601
rect -17 -1743 17 -1709
rect -61 -1969 -27 -1793
rect 27 -1969 61 -1793
rect -17 -2053 17 -2019
rect -17 -2161 17 -2127
rect -61 -2387 -27 -2211
rect 27 -2387 61 -2211
rect -17 -2471 17 -2437
rect -17 -2579 17 -2545
rect -61 -2805 -27 -2629
rect 27 -2805 61 -2629
rect -17 -2889 17 -2855
rect -17 -2997 17 -2963
rect -61 -3223 -27 -3047
rect 27 -3223 61 -3047
rect -17 -3307 17 -3273
rect -17 -3415 17 -3381
rect -61 -3641 -27 -3465
rect 27 -3641 61 -3465
rect -17 -3725 17 -3691
rect -17 -3833 17 -3799
rect -61 -4059 -27 -3883
rect 27 -4059 61 -3883
rect -17 -4143 17 -4109
rect -17 -4251 17 -4217
rect -61 -4477 -27 -4301
rect 27 -4477 61 -4301
rect -17 -4561 17 -4527
rect -17 -4669 17 -4635
rect -61 -4895 -27 -4719
rect 27 -4895 61 -4719
rect -17 -4979 17 -4945
rect -17 -5087 17 -5053
rect -61 -5313 -27 -5137
rect 27 -5313 61 -5137
rect -17 -5397 17 -5363
rect -17 -5505 17 -5471
rect -61 -5731 -27 -5555
rect 27 -5731 61 -5555
rect -17 -5815 17 -5781
<< metal1 >>
rect -29 5815 29 5821
rect -29 5781 -17 5815
rect 17 5781 29 5815
rect -29 5775 29 5781
rect -67 5731 -21 5743
rect -67 5555 -61 5731
rect -27 5555 -21 5731
rect -67 5543 -21 5555
rect 21 5731 67 5743
rect 21 5555 27 5731
rect 61 5555 67 5731
rect 21 5543 67 5555
rect -29 5505 29 5511
rect -29 5471 -17 5505
rect 17 5471 29 5505
rect -29 5465 29 5471
rect -29 5397 29 5403
rect -29 5363 -17 5397
rect 17 5363 29 5397
rect -29 5357 29 5363
rect -67 5313 -21 5325
rect -67 5137 -61 5313
rect -27 5137 -21 5313
rect -67 5125 -21 5137
rect 21 5313 67 5325
rect 21 5137 27 5313
rect 61 5137 67 5313
rect 21 5125 67 5137
rect -29 5087 29 5093
rect -29 5053 -17 5087
rect 17 5053 29 5087
rect -29 5047 29 5053
rect -29 4979 29 4985
rect -29 4945 -17 4979
rect 17 4945 29 4979
rect -29 4939 29 4945
rect -67 4895 -21 4907
rect -67 4719 -61 4895
rect -27 4719 -21 4895
rect -67 4707 -21 4719
rect 21 4895 67 4907
rect 21 4719 27 4895
rect 61 4719 67 4895
rect 21 4707 67 4719
rect -29 4669 29 4675
rect -29 4635 -17 4669
rect 17 4635 29 4669
rect -29 4629 29 4635
rect -29 4561 29 4567
rect -29 4527 -17 4561
rect 17 4527 29 4561
rect -29 4521 29 4527
rect -67 4477 -21 4489
rect -67 4301 -61 4477
rect -27 4301 -21 4477
rect -67 4289 -21 4301
rect 21 4477 67 4489
rect 21 4301 27 4477
rect 61 4301 67 4477
rect 21 4289 67 4301
rect -29 4251 29 4257
rect -29 4217 -17 4251
rect 17 4217 29 4251
rect -29 4211 29 4217
rect -29 4143 29 4149
rect -29 4109 -17 4143
rect 17 4109 29 4143
rect -29 4103 29 4109
rect -67 4059 -21 4071
rect -67 3883 -61 4059
rect -27 3883 -21 4059
rect -67 3871 -21 3883
rect 21 4059 67 4071
rect 21 3883 27 4059
rect 61 3883 67 4059
rect 21 3871 67 3883
rect -29 3833 29 3839
rect -29 3799 -17 3833
rect 17 3799 29 3833
rect -29 3793 29 3799
rect -29 3725 29 3731
rect -29 3691 -17 3725
rect 17 3691 29 3725
rect -29 3685 29 3691
rect -67 3641 -21 3653
rect -67 3465 -61 3641
rect -27 3465 -21 3641
rect -67 3453 -21 3465
rect 21 3641 67 3653
rect 21 3465 27 3641
rect 61 3465 67 3641
rect 21 3453 67 3465
rect -29 3415 29 3421
rect -29 3381 -17 3415
rect 17 3381 29 3415
rect -29 3375 29 3381
rect -29 3307 29 3313
rect -29 3273 -17 3307
rect 17 3273 29 3307
rect -29 3267 29 3273
rect -67 3223 -21 3235
rect -67 3047 -61 3223
rect -27 3047 -21 3223
rect -67 3035 -21 3047
rect 21 3223 67 3235
rect 21 3047 27 3223
rect 61 3047 67 3223
rect 21 3035 67 3047
rect -29 2997 29 3003
rect -29 2963 -17 2997
rect 17 2963 29 2997
rect -29 2957 29 2963
rect -29 2889 29 2895
rect -29 2855 -17 2889
rect 17 2855 29 2889
rect -29 2849 29 2855
rect -67 2805 -21 2817
rect -67 2629 -61 2805
rect -27 2629 -21 2805
rect -67 2617 -21 2629
rect 21 2805 67 2817
rect 21 2629 27 2805
rect 61 2629 67 2805
rect 21 2617 67 2629
rect -29 2579 29 2585
rect -29 2545 -17 2579
rect 17 2545 29 2579
rect -29 2539 29 2545
rect -29 2471 29 2477
rect -29 2437 -17 2471
rect 17 2437 29 2471
rect -29 2431 29 2437
rect -67 2387 -21 2399
rect -67 2211 -61 2387
rect -27 2211 -21 2387
rect -67 2199 -21 2211
rect 21 2387 67 2399
rect 21 2211 27 2387
rect 61 2211 67 2387
rect 21 2199 67 2211
rect -29 2161 29 2167
rect -29 2127 -17 2161
rect 17 2127 29 2161
rect -29 2121 29 2127
rect -29 2053 29 2059
rect -29 2019 -17 2053
rect 17 2019 29 2053
rect -29 2013 29 2019
rect -67 1969 -21 1981
rect -67 1793 -61 1969
rect -27 1793 -21 1969
rect -67 1781 -21 1793
rect 21 1969 67 1981
rect 21 1793 27 1969
rect 61 1793 67 1969
rect 21 1781 67 1793
rect -29 1743 29 1749
rect -29 1709 -17 1743
rect 17 1709 29 1743
rect -29 1703 29 1709
rect -29 1635 29 1641
rect -29 1601 -17 1635
rect 17 1601 29 1635
rect -29 1595 29 1601
rect -67 1551 -21 1563
rect -67 1375 -61 1551
rect -27 1375 -21 1551
rect -67 1363 -21 1375
rect 21 1551 67 1563
rect 21 1375 27 1551
rect 61 1375 67 1551
rect 21 1363 67 1375
rect -29 1325 29 1331
rect -29 1291 -17 1325
rect 17 1291 29 1325
rect -29 1285 29 1291
rect -29 1217 29 1223
rect -29 1183 -17 1217
rect 17 1183 29 1217
rect -29 1177 29 1183
rect -67 1133 -21 1145
rect -67 957 -61 1133
rect -27 957 -21 1133
rect -67 945 -21 957
rect 21 1133 67 1145
rect 21 957 27 1133
rect 61 957 67 1133
rect 21 945 67 957
rect -29 907 29 913
rect -29 873 -17 907
rect 17 873 29 907
rect -29 867 29 873
rect -29 799 29 805
rect -29 765 -17 799
rect 17 765 29 799
rect -29 759 29 765
rect -67 715 -21 727
rect -67 539 -61 715
rect -27 539 -21 715
rect -67 527 -21 539
rect 21 715 67 727
rect 21 539 27 715
rect 61 539 67 715
rect 21 527 67 539
rect -29 489 29 495
rect -29 455 -17 489
rect 17 455 29 489
rect -29 449 29 455
rect -29 381 29 387
rect -29 347 -17 381
rect 17 347 29 381
rect -29 341 29 347
rect -67 297 -21 309
rect -67 121 -61 297
rect -27 121 -21 297
rect -67 109 -21 121
rect 21 297 67 309
rect 21 121 27 297
rect 61 121 67 297
rect 21 109 67 121
rect -29 71 29 77
rect -29 37 -17 71
rect 17 37 29 71
rect -29 31 29 37
rect -29 -37 29 -31
rect -29 -71 -17 -37
rect 17 -71 29 -37
rect -29 -77 29 -71
rect -67 -121 -21 -109
rect -67 -297 -61 -121
rect -27 -297 -21 -121
rect -67 -309 -21 -297
rect 21 -121 67 -109
rect 21 -297 27 -121
rect 61 -297 67 -121
rect 21 -309 67 -297
rect -29 -347 29 -341
rect -29 -381 -17 -347
rect 17 -381 29 -347
rect -29 -387 29 -381
rect -29 -455 29 -449
rect -29 -489 -17 -455
rect 17 -489 29 -455
rect -29 -495 29 -489
rect -67 -539 -21 -527
rect -67 -715 -61 -539
rect -27 -715 -21 -539
rect -67 -727 -21 -715
rect 21 -539 67 -527
rect 21 -715 27 -539
rect 61 -715 67 -539
rect 21 -727 67 -715
rect -29 -765 29 -759
rect -29 -799 -17 -765
rect 17 -799 29 -765
rect -29 -805 29 -799
rect -29 -873 29 -867
rect -29 -907 -17 -873
rect 17 -907 29 -873
rect -29 -913 29 -907
rect -67 -957 -21 -945
rect -67 -1133 -61 -957
rect -27 -1133 -21 -957
rect -67 -1145 -21 -1133
rect 21 -957 67 -945
rect 21 -1133 27 -957
rect 61 -1133 67 -957
rect 21 -1145 67 -1133
rect -29 -1183 29 -1177
rect -29 -1217 -17 -1183
rect 17 -1217 29 -1183
rect -29 -1223 29 -1217
rect -29 -1291 29 -1285
rect -29 -1325 -17 -1291
rect 17 -1325 29 -1291
rect -29 -1331 29 -1325
rect -67 -1375 -21 -1363
rect -67 -1551 -61 -1375
rect -27 -1551 -21 -1375
rect -67 -1563 -21 -1551
rect 21 -1375 67 -1363
rect 21 -1551 27 -1375
rect 61 -1551 67 -1375
rect 21 -1563 67 -1551
rect -29 -1601 29 -1595
rect -29 -1635 -17 -1601
rect 17 -1635 29 -1601
rect -29 -1641 29 -1635
rect -29 -1709 29 -1703
rect -29 -1743 -17 -1709
rect 17 -1743 29 -1709
rect -29 -1749 29 -1743
rect -67 -1793 -21 -1781
rect -67 -1969 -61 -1793
rect -27 -1969 -21 -1793
rect -67 -1981 -21 -1969
rect 21 -1793 67 -1781
rect 21 -1969 27 -1793
rect 61 -1969 67 -1793
rect 21 -1981 67 -1969
rect -29 -2019 29 -2013
rect -29 -2053 -17 -2019
rect 17 -2053 29 -2019
rect -29 -2059 29 -2053
rect -29 -2127 29 -2121
rect -29 -2161 -17 -2127
rect 17 -2161 29 -2127
rect -29 -2167 29 -2161
rect -67 -2211 -21 -2199
rect -67 -2387 -61 -2211
rect -27 -2387 -21 -2211
rect -67 -2399 -21 -2387
rect 21 -2211 67 -2199
rect 21 -2387 27 -2211
rect 61 -2387 67 -2211
rect 21 -2399 67 -2387
rect -29 -2437 29 -2431
rect -29 -2471 -17 -2437
rect 17 -2471 29 -2437
rect -29 -2477 29 -2471
rect -29 -2545 29 -2539
rect -29 -2579 -17 -2545
rect 17 -2579 29 -2545
rect -29 -2585 29 -2579
rect -67 -2629 -21 -2617
rect -67 -2805 -61 -2629
rect -27 -2805 -21 -2629
rect -67 -2817 -21 -2805
rect 21 -2629 67 -2617
rect 21 -2805 27 -2629
rect 61 -2805 67 -2629
rect 21 -2817 67 -2805
rect -29 -2855 29 -2849
rect -29 -2889 -17 -2855
rect 17 -2889 29 -2855
rect -29 -2895 29 -2889
rect -29 -2963 29 -2957
rect -29 -2997 -17 -2963
rect 17 -2997 29 -2963
rect -29 -3003 29 -2997
rect -67 -3047 -21 -3035
rect -67 -3223 -61 -3047
rect -27 -3223 -21 -3047
rect -67 -3235 -21 -3223
rect 21 -3047 67 -3035
rect 21 -3223 27 -3047
rect 61 -3223 67 -3047
rect 21 -3235 67 -3223
rect -29 -3273 29 -3267
rect -29 -3307 -17 -3273
rect 17 -3307 29 -3273
rect -29 -3313 29 -3307
rect -29 -3381 29 -3375
rect -29 -3415 -17 -3381
rect 17 -3415 29 -3381
rect -29 -3421 29 -3415
rect -67 -3465 -21 -3453
rect -67 -3641 -61 -3465
rect -27 -3641 -21 -3465
rect -67 -3653 -21 -3641
rect 21 -3465 67 -3453
rect 21 -3641 27 -3465
rect 61 -3641 67 -3465
rect 21 -3653 67 -3641
rect -29 -3691 29 -3685
rect -29 -3725 -17 -3691
rect 17 -3725 29 -3691
rect -29 -3731 29 -3725
rect -29 -3799 29 -3793
rect -29 -3833 -17 -3799
rect 17 -3833 29 -3799
rect -29 -3839 29 -3833
rect -67 -3883 -21 -3871
rect -67 -4059 -61 -3883
rect -27 -4059 -21 -3883
rect -67 -4071 -21 -4059
rect 21 -3883 67 -3871
rect 21 -4059 27 -3883
rect 61 -4059 67 -3883
rect 21 -4071 67 -4059
rect -29 -4109 29 -4103
rect -29 -4143 -17 -4109
rect 17 -4143 29 -4109
rect -29 -4149 29 -4143
rect -29 -4217 29 -4211
rect -29 -4251 -17 -4217
rect 17 -4251 29 -4217
rect -29 -4257 29 -4251
rect -67 -4301 -21 -4289
rect -67 -4477 -61 -4301
rect -27 -4477 -21 -4301
rect -67 -4489 -21 -4477
rect 21 -4301 67 -4289
rect 21 -4477 27 -4301
rect 61 -4477 67 -4301
rect 21 -4489 67 -4477
rect -29 -4527 29 -4521
rect -29 -4561 -17 -4527
rect 17 -4561 29 -4527
rect -29 -4567 29 -4561
rect -29 -4635 29 -4629
rect -29 -4669 -17 -4635
rect 17 -4669 29 -4635
rect -29 -4675 29 -4669
rect -67 -4719 -21 -4707
rect -67 -4895 -61 -4719
rect -27 -4895 -21 -4719
rect -67 -4907 -21 -4895
rect 21 -4719 67 -4707
rect 21 -4895 27 -4719
rect 61 -4895 67 -4719
rect 21 -4907 67 -4895
rect -29 -4945 29 -4939
rect -29 -4979 -17 -4945
rect 17 -4979 29 -4945
rect -29 -4985 29 -4979
rect -29 -5053 29 -5047
rect -29 -5087 -17 -5053
rect 17 -5087 29 -5053
rect -29 -5093 29 -5087
rect -67 -5137 -21 -5125
rect -67 -5313 -61 -5137
rect -27 -5313 -21 -5137
rect -67 -5325 -21 -5313
rect 21 -5137 67 -5125
rect 21 -5313 27 -5137
rect 61 -5313 67 -5137
rect 21 -5325 67 -5313
rect -29 -5363 29 -5357
rect -29 -5397 -17 -5363
rect 17 -5397 29 -5363
rect -29 -5403 29 -5397
rect -29 -5471 29 -5465
rect -29 -5505 -17 -5471
rect 17 -5505 29 -5471
rect -29 -5511 29 -5505
rect -67 -5555 -21 -5543
rect -67 -5731 -61 -5555
rect -27 -5731 -21 -5555
rect -67 -5743 -21 -5731
rect 21 -5555 67 -5543
rect 21 -5731 27 -5555
rect 61 -5731 67 -5555
rect 21 -5743 67 -5731
rect -29 -5781 29 -5775
rect -29 -5815 -17 -5781
rect 17 -5815 29 -5781
rect -29 -5821 29 -5815
<< properties >>
string FIXED_BBOX -158 -5900 158 5900
string gencell sky130_fd_pr__nfet_01v8_lvt
string library sky130
string parameters w 1 l 0.150 m 28 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
