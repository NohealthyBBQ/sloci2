magic
tech sky130A
magscale 1 2
timestamp 1662302892
<< pwell >>
rect -625 -1646 625 1646
<< nmoslvt >>
rect -429 1036 -29 1436
rect 29 1036 429 1436
rect -429 418 -29 818
rect 29 418 429 818
rect -429 -200 -29 200
rect 29 -200 429 200
rect -429 -818 -29 -418
rect 29 -818 429 -418
rect -429 -1436 -29 -1036
rect 29 -1436 429 -1036
<< ndiff >>
rect -487 1424 -429 1436
rect -487 1048 -475 1424
rect -441 1048 -429 1424
rect -487 1036 -429 1048
rect -29 1424 29 1436
rect -29 1048 -17 1424
rect 17 1048 29 1424
rect -29 1036 29 1048
rect 429 1424 487 1436
rect 429 1048 441 1424
rect 475 1048 487 1424
rect 429 1036 487 1048
rect -487 806 -429 818
rect -487 430 -475 806
rect -441 430 -429 806
rect -487 418 -429 430
rect -29 806 29 818
rect -29 430 -17 806
rect 17 430 29 806
rect -29 418 29 430
rect 429 806 487 818
rect 429 430 441 806
rect 475 430 487 806
rect 429 418 487 430
rect -487 188 -429 200
rect -487 -188 -475 188
rect -441 -188 -429 188
rect -487 -200 -429 -188
rect -29 188 29 200
rect -29 -188 -17 188
rect 17 -188 29 188
rect -29 -200 29 -188
rect 429 188 487 200
rect 429 -188 441 188
rect 475 -188 487 188
rect 429 -200 487 -188
rect -487 -430 -429 -418
rect -487 -806 -475 -430
rect -441 -806 -429 -430
rect -487 -818 -429 -806
rect -29 -430 29 -418
rect -29 -806 -17 -430
rect 17 -806 29 -430
rect -29 -818 29 -806
rect 429 -430 487 -418
rect 429 -806 441 -430
rect 475 -806 487 -430
rect 429 -818 487 -806
rect -487 -1048 -429 -1036
rect -487 -1424 -475 -1048
rect -441 -1424 -429 -1048
rect -487 -1436 -429 -1424
rect -29 -1048 29 -1036
rect -29 -1424 -17 -1048
rect 17 -1424 29 -1048
rect -29 -1436 29 -1424
rect 429 -1048 487 -1036
rect 429 -1424 441 -1048
rect 475 -1424 487 -1048
rect 429 -1436 487 -1424
<< ndiffc >>
rect -475 1048 -441 1424
rect -17 1048 17 1424
rect 441 1048 475 1424
rect -475 430 -441 806
rect -17 430 17 806
rect 441 430 475 806
rect -475 -188 -441 188
rect -17 -188 17 188
rect 441 -188 475 188
rect -475 -806 -441 -430
rect -17 -806 17 -430
rect 441 -806 475 -430
rect -475 -1424 -441 -1048
rect -17 -1424 17 -1048
rect 441 -1424 475 -1048
<< psubdiff >>
rect -589 1576 -493 1610
rect 493 1576 589 1610
rect -589 1514 -555 1576
rect 555 1514 589 1576
rect -589 -1576 -555 -1514
rect 555 -1576 589 -1514
rect -589 -1610 -493 -1576
rect 493 -1610 589 -1576
<< psubdiffcont >>
rect -493 1576 493 1610
rect -589 -1514 -555 1514
rect 555 -1514 589 1514
rect -493 -1610 493 -1576
<< poly >>
rect -429 1508 -29 1524
rect -429 1474 -413 1508
rect -45 1474 -29 1508
rect -429 1436 -29 1474
rect 29 1508 429 1524
rect 29 1474 45 1508
rect 413 1474 429 1508
rect 29 1436 429 1474
rect -429 998 -29 1036
rect -429 964 -413 998
rect -45 964 -29 998
rect -429 948 -29 964
rect 29 998 429 1036
rect 29 964 45 998
rect 413 964 429 998
rect 29 948 429 964
rect -429 890 -29 906
rect -429 856 -413 890
rect -45 856 -29 890
rect -429 818 -29 856
rect 29 890 429 906
rect 29 856 45 890
rect 413 856 429 890
rect 29 818 429 856
rect -429 380 -29 418
rect -429 346 -413 380
rect -45 346 -29 380
rect -429 330 -29 346
rect 29 380 429 418
rect 29 346 45 380
rect 413 346 429 380
rect 29 330 429 346
rect -429 272 -29 288
rect -429 238 -413 272
rect -45 238 -29 272
rect -429 200 -29 238
rect 29 272 429 288
rect 29 238 45 272
rect 413 238 429 272
rect 29 200 429 238
rect -429 -238 -29 -200
rect -429 -272 -413 -238
rect -45 -272 -29 -238
rect -429 -288 -29 -272
rect 29 -238 429 -200
rect 29 -272 45 -238
rect 413 -272 429 -238
rect 29 -288 429 -272
rect -429 -346 -29 -330
rect -429 -380 -413 -346
rect -45 -380 -29 -346
rect -429 -418 -29 -380
rect 29 -346 429 -330
rect 29 -380 45 -346
rect 413 -380 429 -346
rect 29 -418 429 -380
rect -429 -856 -29 -818
rect -429 -890 -413 -856
rect -45 -890 -29 -856
rect -429 -906 -29 -890
rect 29 -856 429 -818
rect 29 -890 45 -856
rect 413 -890 429 -856
rect 29 -906 429 -890
rect -429 -964 -29 -948
rect -429 -998 -413 -964
rect -45 -998 -29 -964
rect -429 -1036 -29 -998
rect 29 -964 429 -948
rect 29 -998 45 -964
rect 413 -998 429 -964
rect 29 -1036 429 -998
rect -429 -1474 -29 -1436
rect -429 -1508 -413 -1474
rect -45 -1508 -29 -1474
rect -429 -1524 -29 -1508
rect 29 -1474 429 -1436
rect 29 -1508 45 -1474
rect 413 -1508 429 -1474
rect 29 -1524 429 -1508
<< polycont >>
rect -413 1474 -45 1508
rect 45 1474 413 1508
rect -413 964 -45 998
rect 45 964 413 998
rect -413 856 -45 890
rect 45 856 413 890
rect -413 346 -45 380
rect 45 346 413 380
rect -413 238 -45 272
rect 45 238 413 272
rect -413 -272 -45 -238
rect 45 -272 413 -238
rect -413 -380 -45 -346
rect 45 -380 413 -346
rect -413 -890 -45 -856
rect 45 -890 413 -856
rect -413 -998 -45 -964
rect 45 -998 413 -964
rect -413 -1508 -45 -1474
rect 45 -1508 413 -1474
<< locali >>
rect -589 1576 -493 1610
rect 493 1576 589 1610
rect -589 1514 -555 1576
rect 555 1514 589 1576
rect -429 1474 -413 1508
rect -45 1474 -29 1508
rect 29 1474 45 1508
rect 413 1474 429 1508
rect -475 1424 -441 1440
rect -475 1032 -441 1048
rect -17 1424 17 1440
rect -17 1032 17 1048
rect 441 1424 475 1440
rect 441 1032 475 1048
rect -429 964 -413 998
rect -45 964 -29 998
rect 29 964 45 998
rect 413 964 429 998
rect -429 856 -413 890
rect -45 856 -29 890
rect 29 856 45 890
rect 413 856 429 890
rect -475 806 -441 822
rect -475 414 -441 430
rect -17 806 17 822
rect -17 414 17 430
rect 441 806 475 822
rect 441 414 475 430
rect -429 346 -413 380
rect -45 346 -29 380
rect 29 346 45 380
rect 413 346 429 380
rect -429 238 -413 272
rect -45 238 -29 272
rect 29 238 45 272
rect 413 238 429 272
rect -475 188 -441 204
rect -475 -204 -441 -188
rect -17 188 17 204
rect -17 -204 17 -188
rect 441 188 475 204
rect 441 -204 475 -188
rect -429 -272 -413 -238
rect -45 -272 -29 -238
rect 29 -272 45 -238
rect 413 -272 429 -238
rect -429 -380 -413 -346
rect -45 -380 -29 -346
rect 29 -380 45 -346
rect 413 -380 429 -346
rect -475 -430 -441 -414
rect -475 -822 -441 -806
rect -17 -430 17 -414
rect -17 -822 17 -806
rect 441 -430 475 -414
rect 441 -822 475 -806
rect -429 -890 -413 -856
rect -45 -890 -29 -856
rect 29 -890 45 -856
rect 413 -890 429 -856
rect -429 -998 -413 -964
rect -45 -998 -29 -964
rect 29 -998 45 -964
rect 413 -998 429 -964
rect -475 -1048 -441 -1032
rect -475 -1440 -441 -1424
rect -17 -1048 17 -1032
rect -17 -1440 17 -1424
rect 441 -1048 475 -1032
rect 441 -1440 475 -1424
rect -429 -1508 -413 -1474
rect -45 -1508 -29 -1474
rect 29 -1508 45 -1474
rect 413 -1508 429 -1474
rect -589 -1576 -555 -1514
rect 555 -1576 589 -1514
rect -589 -1610 -493 -1576
rect 493 -1610 589 -1576
<< viali >>
rect -413 1474 -45 1508
rect 45 1474 413 1508
rect -475 1048 -441 1424
rect -17 1048 17 1424
rect 441 1048 475 1424
rect -413 964 -45 998
rect 45 964 413 998
rect -413 856 -45 890
rect 45 856 413 890
rect -475 430 -441 806
rect -17 430 17 806
rect 441 430 475 806
rect -413 346 -45 380
rect 45 346 413 380
rect -413 238 -45 272
rect 45 238 413 272
rect -475 -188 -441 188
rect -17 -188 17 188
rect 441 -188 475 188
rect -413 -272 -45 -238
rect 45 -272 413 -238
rect -413 -380 -45 -346
rect 45 -380 413 -346
rect -475 -806 -441 -430
rect -17 -806 17 -430
rect 441 -806 475 -430
rect -413 -890 -45 -856
rect 45 -890 413 -856
rect -413 -998 -45 -964
rect 45 -998 413 -964
rect -475 -1424 -441 -1048
rect -17 -1424 17 -1048
rect 441 -1424 475 -1048
rect -413 -1508 -45 -1474
rect 45 -1508 413 -1474
<< metal1 >>
rect -425 1508 -33 1514
rect -425 1474 -413 1508
rect -45 1474 -33 1508
rect -425 1468 -33 1474
rect 33 1508 425 1514
rect 33 1474 45 1508
rect 413 1474 425 1508
rect 33 1468 425 1474
rect -481 1424 -435 1436
rect -481 1048 -475 1424
rect -441 1048 -435 1424
rect -481 1036 -435 1048
rect -23 1424 23 1436
rect -23 1048 -17 1424
rect 17 1048 23 1424
rect -23 1036 23 1048
rect 435 1424 481 1436
rect 435 1048 441 1424
rect 475 1048 481 1424
rect 435 1036 481 1048
rect -425 998 -33 1004
rect -425 964 -413 998
rect -45 964 -33 998
rect -425 958 -33 964
rect 33 998 425 1004
rect 33 964 45 998
rect 413 964 425 998
rect 33 958 425 964
rect -425 890 -33 896
rect -425 856 -413 890
rect -45 856 -33 890
rect -425 850 -33 856
rect 33 890 425 896
rect 33 856 45 890
rect 413 856 425 890
rect 33 850 425 856
rect -481 806 -435 818
rect -481 430 -475 806
rect -441 430 -435 806
rect -481 418 -435 430
rect -23 806 23 818
rect -23 430 -17 806
rect 17 430 23 806
rect -23 418 23 430
rect 435 806 481 818
rect 435 430 441 806
rect 475 430 481 806
rect 435 418 481 430
rect -425 380 -33 386
rect -425 346 -413 380
rect -45 346 -33 380
rect -425 340 -33 346
rect 33 380 425 386
rect 33 346 45 380
rect 413 346 425 380
rect 33 340 425 346
rect -425 272 -33 278
rect -425 238 -413 272
rect -45 238 -33 272
rect -425 232 -33 238
rect 33 272 425 278
rect 33 238 45 272
rect 413 238 425 272
rect 33 232 425 238
rect -481 188 -435 200
rect -481 -188 -475 188
rect -441 -188 -435 188
rect -481 -200 -435 -188
rect -23 188 23 200
rect -23 -188 -17 188
rect 17 -188 23 188
rect -23 -200 23 -188
rect 435 188 481 200
rect 435 -188 441 188
rect 475 -188 481 188
rect 435 -200 481 -188
rect -425 -238 -33 -232
rect -425 -272 -413 -238
rect -45 -272 -33 -238
rect -425 -278 -33 -272
rect 33 -238 425 -232
rect 33 -272 45 -238
rect 413 -272 425 -238
rect 33 -278 425 -272
rect -425 -346 -33 -340
rect -425 -380 -413 -346
rect -45 -380 -33 -346
rect -425 -386 -33 -380
rect 33 -346 425 -340
rect 33 -380 45 -346
rect 413 -380 425 -346
rect 33 -386 425 -380
rect -481 -430 -435 -418
rect -481 -806 -475 -430
rect -441 -806 -435 -430
rect -481 -818 -435 -806
rect -23 -430 23 -418
rect -23 -806 -17 -430
rect 17 -806 23 -430
rect -23 -818 23 -806
rect 435 -430 481 -418
rect 435 -806 441 -430
rect 475 -806 481 -430
rect 435 -818 481 -806
rect -425 -856 -33 -850
rect -425 -890 -413 -856
rect -45 -890 -33 -856
rect -425 -896 -33 -890
rect 33 -856 425 -850
rect 33 -890 45 -856
rect 413 -890 425 -856
rect 33 -896 425 -890
rect -425 -964 -33 -958
rect -425 -998 -413 -964
rect -45 -998 -33 -964
rect -425 -1004 -33 -998
rect 33 -964 425 -958
rect 33 -998 45 -964
rect 413 -998 425 -964
rect 33 -1004 425 -998
rect -481 -1048 -435 -1036
rect -481 -1424 -475 -1048
rect -441 -1424 -435 -1048
rect -481 -1436 -435 -1424
rect -23 -1048 23 -1036
rect -23 -1424 -17 -1048
rect 17 -1424 23 -1048
rect -23 -1436 23 -1424
rect 435 -1048 481 -1036
rect 435 -1424 441 -1048
rect 475 -1424 481 -1048
rect 435 -1436 481 -1424
rect -425 -1474 -33 -1468
rect -425 -1508 -413 -1474
rect -45 -1508 -33 -1474
rect -425 -1514 -33 -1508
rect 33 -1474 425 -1468
rect 33 -1508 45 -1474
rect 413 -1508 425 -1474
rect 33 -1514 425 -1508
<< properties >>
string FIXED_BBOX -572 -1593 572 1593
string gencell sky130_fd_pr__nfet_01v8_lvt
string library sky130
string parameters w 2 l 2 m 5 nf 2 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
