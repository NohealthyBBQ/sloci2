magic
tech sky130A
magscale 1 2
timestamp 1671759029
<< nwell >>
rect -1999 -1819 1999 1819
<< pmoslvt >>
rect -1803 -1600 -1403 1600
rect -1345 -1600 -945 1600
rect -887 -1600 -487 1600
rect -429 -1600 -29 1600
rect 29 -1600 429 1600
rect 487 -1600 887 1600
rect 945 -1600 1345 1600
rect 1403 -1600 1803 1600
<< pdiff >>
rect -1861 1588 -1803 1600
rect -1861 -1588 -1849 1588
rect -1815 -1588 -1803 1588
rect -1861 -1600 -1803 -1588
rect -1403 1588 -1345 1600
rect -1403 -1588 -1391 1588
rect -1357 -1588 -1345 1588
rect -1403 -1600 -1345 -1588
rect -945 1588 -887 1600
rect -945 -1588 -933 1588
rect -899 -1588 -887 1588
rect -945 -1600 -887 -1588
rect -487 1588 -429 1600
rect -487 -1588 -475 1588
rect -441 -1588 -429 1588
rect -487 -1600 -429 -1588
rect -29 1588 29 1600
rect -29 -1588 -17 1588
rect 17 -1588 29 1588
rect -29 -1600 29 -1588
rect 429 1588 487 1600
rect 429 -1588 441 1588
rect 475 -1588 487 1588
rect 429 -1600 487 -1588
rect 887 1588 945 1600
rect 887 -1588 899 1588
rect 933 -1588 945 1588
rect 887 -1600 945 -1588
rect 1345 1588 1403 1600
rect 1345 -1588 1357 1588
rect 1391 -1588 1403 1588
rect 1345 -1600 1403 -1588
rect 1803 1588 1861 1600
rect 1803 -1588 1815 1588
rect 1849 -1588 1861 1588
rect 1803 -1600 1861 -1588
<< pdiffc >>
rect -1849 -1588 -1815 1588
rect -1391 -1588 -1357 1588
rect -933 -1588 -899 1588
rect -475 -1588 -441 1588
rect -17 -1588 17 1588
rect 441 -1588 475 1588
rect 899 -1588 933 1588
rect 1357 -1588 1391 1588
rect 1815 -1588 1849 1588
<< nsubdiff >>
rect -1963 1749 -1867 1783
rect 1867 1749 1963 1783
rect -1963 1687 -1929 1749
rect 1929 1687 1963 1749
rect -1963 -1749 -1929 -1687
rect 1929 -1749 1963 -1687
rect -1963 -1783 -1867 -1749
rect 1867 -1783 1963 -1749
<< nsubdiffcont >>
rect -1867 1749 1867 1783
rect -1963 -1687 -1929 1687
rect 1929 -1687 1963 1687
rect -1867 -1783 1867 -1749
<< poly >>
rect -1803 1681 -1403 1697
rect -1803 1647 -1787 1681
rect -1419 1647 -1403 1681
rect -1803 1600 -1403 1647
rect -1345 1681 -945 1697
rect -1345 1647 -1329 1681
rect -961 1647 -945 1681
rect -1345 1600 -945 1647
rect -887 1681 -487 1697
rect -887 1647 -871 1681
rect -503 1647 -487 1681
rect -887 1600 -487 1647
rect -429 1681 -29 1697
rect -429 1647 -413 1681
rect -45 1647 -29 1681
rect -429 1600 -29 1647
rect 29 1681 429 1697
rect 29 1647 45 1681
rect 413 1647 429 1681
rect 29 1600 429 1647
rect 487 1681 887 1697
rect 487 1647 503 1681
rect 871 1647 887 1681
rect 487 1600 887 1647
rect 945 1681 1345 1697
rect 945 1647 961 1681
rect 1329 1647 1345 1681
rect 945 1600 1345 1647
rect 1403 1681 1803 1697
rect 1403 1647 1419 1681
rect 1787 1647 1803 1681
rect 1403 1600 1803 1647
rect -1803 -1647 -1403 -1600
rect -1803 -1681 -1787 -1647
rect -1419 -1681 -1403 -1647
rect -1803 -1697 -1403 -1681
rect -1345 -1647 -945 -1600
rect -1345 -1681 -1329 -1647
rect -961 -1681 -945 -1647
rect -1345 -1697 -945 -1681
rect -887 -1647 -487 -1600
rect -887 -1681 -871 -1647
rect -503 -1681 -487 -1647
rect -887 -1697 -487 -1681
rect -429 -1647 -29 -1600
rect -429 -1681 -413 -1647
rect -45 -1681 -29 -1647
rect -429 -1697 -29 -1681
rect 29 -1647 429 -1600
rect 29 -1681 45 -1647
rect 413 -1681 429 -1647
rect 29 -1697 429 -1681
rect 487 -1647 887 -1600
rect 487 -1681 503 -1647
rect 871 -1681 887 -1647
rect 487 -1697 887 -1681
rect 945 -1647 1345 -1600
rect 945 -1681 961 -1647
rect 1329 -1681 1345 -1647
rect 945 -1697 1345 -1681
rect 1403 -1647 1803 -1600
rect 1403 -1681 1419 -1647
rect 1787 -1681 1803 -1647
rect 1403 -1697 1803 -1681
<< polycont >>
rect -1787 1647 -1419 1681
rect -1329 1647 -961 1681
rect -871 1647 -503 1681
rect -413 1647 -45 1681
rect 45 1647 413 1681
rect 503 1647 871 1681
rect 961 1647 1329 1681
rect 1419 1647 1787 1681
rect -1787 -1681 -1419 -1647
rect -1329 -1681 -961 -1647
rect -871 -1681 -503 -1647
rect -413 -1681 -45 -1647
rect 45 -1681 413 -1647
rect 503 -1681 871 -1647
rect 961 -1681 1329 -1647
rect 1419 -1681 1787 -1647
<< locali >>
rect -1963 1749 -1867 1783
rect 1867 1749 1963 1783
rect -1963 1687 -1929 1749
rect 1929 1687 1963 1749
rect -1803 1647 -1787 1681
rect -1419 1647 -1403 1681
rect -1345 1647 -1329 1681
rect -961 1647 -945 1681
rect -887 1647 -871 1681
rect -503 1647 -487 1681
rect -429 1647 -413 1681
rect -45 1647 -29 1681
rect 29 1647 45 1681
rect 413 1647 429 1681
rect 487 1647 503 1681
rect 871 1647 887 1681
rect 945 1647 961 1681
rect 1329 1647 1345 1681
rect 1403 1647 1419 1681
rect 1787 1647 1803 1681
rect -1849 1588 -1815 1604
rect -1849 -1604 -1815 -1588
rect -1391 1588 -1357 1604
rect -1391 -1604 -1357 -1588
rect -933 1588 -899 1604
rect -933 -1604 -899 -1588
rect -475 1588 -441 1604
rect -475 -1604 -441 -1588
rect -17 1588 17 1604
rect -17 -1604 17 -1588
rect 441 1588 475 1604
rect 441 -1604 475 -1588
rect 899 1588 933 1604
rect 899 -1604 933 -1588
rect 1357 1588 1391 1604
rect 1357 -1604 1391 -1588
rect 1815 1588 1849 1604
rect 1815 -1604 1849 -1588
rect -1803 -1681 -1787 -1647
rect -1419 -1681 -1403 -1647
rect -1345 -1681 -1329 -1647
rect -961 -1681 -945 -1647
rect -887 -1681 -871 -1647
rect -503 -1681 -487 -1647
rect -429 -1681 -413 -1647
rect -45 -1681 -29 -1647
rect 29 -1681 45 -1647
rect 413 -1681 429 -1647
rect 487 -1681 503 -1647
rect 871 -1681 887 -1647
rect 945 -1681 961 -1647
rect 1329 -1681 1345 -1647
rect 1403 -1681 1419 -1647
rect 1787 -1681 1803 -1647
rect -1963 -1749 -1929 -1687
rect 1929 -1749 1963 -1687
rect -1963 -1783 -1867 -1749
rect 1867 -1783 1963 -1749
<< viali >>
rect -1787 1647 -1419 1681
rect -1329 1647 -961 1681
rect -871 1647 -503 1681
rect -413 1647 -45 1681
rect 45 1647 413 1681
rect 503 1647 871 1681
rect 961 1647 1329 1681
rect 1419 1647 1787 1681
rect -1849 -1588 -1815 1588
rect -1391 -1588 -1357 1588
rect -933 -1588 -899 1588
rect -475 -1588 -441 1588
rect -17 -1588 17 1588
rect 441 -1588 475 1588
rect 899 -1588 933 1588
rect 1357 -1588 1391 1588
rect 1815 -1588 1849 1588
rect -1787 -1681 -1419 -1647
rect -1329 -1681 -961 -1647
rect -871 -1681 -503 -1647
rect -413 -1681 -45 -1647
rect 45 -1681 413 -1647
rect 503 -1681 871 -1647
rect 961 -1681 1329 -1647
rect 1419 -1681 1787 -1647
<< metal1 >>
rect -1799 1681 -1407 1687
rect -1799 1647 -1787 1681
rect -1419 1647 -1407 1681
rect -1799 1641 -1407 1647
rect -1341 1681 -949 1687
rect -1341 1647 -1329 1681
rect -961 1647 -949 1681
rect -1341 1641 -949 1647
rect -883 1681 -491 1687
rect -883 1647 -871 1681
rect -503 1647 -491 1681
rect -883 1641 -491 1647
rect -425 1681 -33 1687
rect -425 1647 -413 1681
rect -45 1647 -33 1681
rect -425 1641 -33 1647
rect 33 1681 425 1687
rect 33 1647 45 1681
rect 413 1647 425 1681
rect 33 1641 425 1647
rect 491 1681 883 1687
rect 491 1647 503 1681
rect 871 1647 883 1681
rect 491 1641 883 1647
rect 949 1681 1341 1687
rect 949 1647 961 1681
rect 1329 1647 1341 1681
rect 949 1641 1341 1647
rect 1407 1681 1799 1687
rect 1407 1647 1419 1681
rect 1787 1647 1799 1681
rect 1407 1641 1799 1647
rect -1855 1588 -1809 1600
rect -1855 -1588 -1849 1588
rect -1815 -1588 -1809 1588
rect -1855 -1600 -1809 -1588
rect -1397 1588 -1351 1600
rect -1397 -1588 -1391 1588
rect -1357 -1588 -1351 1588
rect -1397 -1600 -1351 -1588
rect -939 1588 -893 1600
rect -939 -1588 -933 1588
rect -899 -1588 -893 1588
rect -939 -1600 -893 -1588
rect -481 1588 -435 1600
rect -481 -1588 -475 1588
rect -441 -1588 -435 1588
rect -481 -1600 -435 -1588
rect -23 1588 23 1600
rect -23 -1588 -17 1588
rect 17 -1588 23 1588
rect -23 -1600 23 -1588
rect 435 1588 481 1600
rect 435 -1588 441 1588
rect 475 -1588 481 1588
rect 435 -1600 481 -1588
rect 893 1588 939 1600
rect 893 -1588 899 1588
rect 933 -1588 939 1588
rect 893 -1600 939 -1588
rect 1351 1588 1397 1600
rect 1351 -1588 1357 1588
rect 1391 -1588 1397 1588
rect 1351 -1600 1397 -1588
rect 1809 1588 1855 1600
rect 1809 -1588 1815 1588
rect 1849 -1588 1855 1588
rect 1809 -1600 1855 -1588
rect -1799 -1647 -1407 -1641
rect -1799 -1681 -1787 -1647
rect -1419 -1681 -1407 -1647
rect -1799 -1687 -1407 -1681
rect -1341 -1647 -949 -1641
rect -1341 -1681 -1329 -1647
rect -961 -1681 -949 -1647
rect -1341 -1687 -949 -1681
rect -883 -1647 -491 -1641
rect -883 -1681 -871 -1647
rect -503 -1681 -491 -1647
rect -883 -1687 -491 -1681
rect -425 -1647 -33 -1641
rect -425 -1681 -413 -1647
rect -45 -1681 -33 -1647
rect -425 -1687 -33 -1681
rect 33 -1647 425 -1641
rect 33 -1681 45 -1647
rect 413 -1681 425 -1647
rect 33 -1687 425 -1681
rect 491 -1647 883 -1641
rect 491 -1681 503 -1647
rect 871 -1681 883 -1647
rect 491 -1687 883 -1681
rect 949 -1647 1341 -1641
rect 949 -1681 961 -1647
rect 1329 -1681 1341 -1647
rect 949 -1687 1341 -1681
rect 1407 -1647 1799 -1641
rect 1407 -1681 1419 -1647
rect 1787 -1681 1799 -1647
rect 1407 -1687 1799 -1681
<< properties >>
string FIXED_BBOX -1946 -1766 1946 1766
string gencell sky130_fd_pr__pfet_01v8_lvt
string library sky130
string parameters w 16 l 2 m 1 nf 8 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.35 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
