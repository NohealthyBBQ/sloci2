magic
tech sky130A
timestamp 1671754915
<< pwell >>
rect -324 -155 323 155
<< nmoslvt >>
rect -224 -50 -209 50
rect -176 -50 -161 50
rect -128 -50 -113 50
rect -80 -50 -65 50
rect -32 -50 -17 50
rect 16 -50 31 50
rect 64 -50 79 50
rect 112 -50 127 50
rect 160 -50 175 50
rect 208 -50 223 50
<< ndiff >>
rect -255 44 -224 50
rect -255 -44 -249 44
rect -232 -44 -224 44
rect -255 -50 -224 -44
rect -209 44 -176 50
rect -209 -44 -201 44
rect -184 -44 -176 44
rect -209 -50 -176 -44
rect -161 44 -128 50
rect -161 -44 -153 44
rect -136 -44 -128 44
rect -161 -50 -128 -44
rect -113 44 -80 50
rect -113 -44 -105 44
rect -88 -44 -80 44
rect -113 -50 -80 -44
rect -65 44 -32 50
rect -65 -44 -57 44
rect -40 -44 -32 44
rect -65 -50 -32 -44
rect -17 44 16 50
rect -17 -44 -9 44
rect 8 -44 16 44
rect -17 -50 16 -44
rect 31 44 64 50
rect 31 -44 39 44
rect 56 -44 64 44
rect 31 -50 64 -44
rect 79 44 112 50
rect 79 -44 87 44
rect 104 -44 112 44
rect 79 -50 112 -44
rect 127 44 160 50
rect 127 -44 135 44
rect 152 -44 160 44
rect 127 -50 160 -44
rect 175 44 208 50
rect 175 -44 183 44
rect 200 -44 208 44
rect 175 -50 208 -44
rect 223 44 254 50
rect 223 -44 231 44
rect 248 -44 254 44
rect 223 -50 254 -44
<< ndiffc >>
rect -249 -44 -232 44
rect -201 -44 -184 44
rect -153 -44 -136 44
rect -105 -44 -88 44
rect -57 -44 -40 44
rect -9 -44 8 44
rect 39 -44 56 44
rect 87 -44 104 44
rect 135 -44 152 44
rect 183 -44 200 44
rect 231 -44 248 44
<< psubdiff >>
rect -306 120 -258 137
rect 257 120 305 137
rect -306 89 -289 120
rect 288 89 305 120
rect -306 -120 -289 -89
rect 288 -120 305 -89
rect -306 -137 -258 -120
rect 257 -137 305 -120
<< psubdiffcont >>
rect -258 120 257 137
rect -306 -89 -289 89
rect 288 -89 305 89
rect -258 -137 257 -120
<< poly >>
rect -224 50 -209 63
rect -176 50 -161 63
rect -128 50 -113 63
rect -80 50 -65 63
rect -32 50 -17 63
rect 16 50 31 63
rect 64 50 79 63
rect 112 50 127 63
rect 160 50 175 63
rect 208 50 223 63
rect -224 -61 -209 -50
rect -233 -69 -200 -61
rect -176 -69 -161 -50
rect -128 -61 -113 -50
rect -137 -69 -104 -61
rect -80 -69 -65 -50
rect -32 -61 -17 -50
rect -41 -69 -8 -61
rect 16 -69 31 -50
rect 64 -61 79 -50
rect 55 -69 88 -61
rect 112 -69 127 -50
rect 160 -61 175 -50
rect 151 -69 184 -61
rect 208 -69 223 -50
rect -233 -86 -33 -69
rect -16 -86 223 -69
rect -233 -89 223 -86
rect -233 -94 -200 -89
rect -137 -94 -104 -89
rect -41 -94 -8 -89
rect 55 -94 88 -89
rect 151 -94 184 -89
<< polycont >>
rect -33 -86 -16 -69
<< locali >>
rect -306 120 -258 137
rect 257 120 305 137
rect -306 89 -289 120
rect 288 89 305 120
rect -249 44 -232 52
rect -249 -52 -232 -44
rect -201 44 -184 52
rect -201 -52 -184 -44
rect -153 44 -136 52
rect -153 -52 -136 -44
rect -105 44 -88 52
rect -105 -52 -88 -44
rect -57 44 -40 52
rect -57 -52 -40 -44
rect -9 44 8 52
rect -9 -52 8 -44
rect 39 44 56 52
rect 39 -52 56 -44
rect 87 44 104 52
rect 87 -52 104 -44
rect 135 44 152 52
rect 135 -52 152 -44
rect 183 44 200 52
rect 183 -52 200 -44
rect 231 44 248 52
rect 231 -52 248 -44
rect -41 -86 -33 -69
rect -16 -86 -8 -69
rect -306 -120 -289 -89
rect 288 -120 305 -89
rect -306 -137 -258 -120
rect 257 -137 305 -120
<< viali >>
rect -249 -44 -232 44
rect -201 -44 -184 44
rect -153 -44 -136 44
rect -105 -44 -88 44
rect -57 -44 -40 44
rect -9 -44 8 44
rect 39 -44 56 44
rect 87 -44 104 44
rect 135 -44 152 44
rect 183 -44 200 44
rect 231 -44 248 44
rect -33 -86 -16 -69
<< metal1 >>
rect -252 44 -229 50
rect -252 -15 -249 44
rect -257 -18 -249 -15
rect -232 -15 -229 44
rect -209 48 -176 50
rect -209 18 -205 48
rect -179 18 -176 48
rect -209 15 -201 18
rect -232 -18 -224 -15
rect -257 -48 -254 -18
rect -228 -48 -224 -18
rect -257 -50 -224 -48
rect -204 -44 -201 15
rect -184 15 -176 18
rect -156 44 -133 50
rect -184 -44 -181 15
rect -156 -15 -153 44
rect -204 -50 -181 -44
rect -161 -17 -153 -15
rect -136 -15 -133 44
rect -113 48 -80 50
rect -113 18 -109 48
rect -83 18 -80 48
rect -113 15 -105 18
rect -136 -17 -128 -15
rect -161 -47 -157 -17
rect -131 -47 -128 -17
rect -161 -50 -128 -47
rect -108 -44 -105 15
rect -88 15 -80 18
rect -60 44 -37 50
rect -88 -44 -85 15
rect -60 -15 -57 44
rect -108 -50 -85 -44
rect -65 -17 -57 -15
rect -40 -15 -37 44
rect -17 48 16 50
rect -17 18 -14 48
rect 12 18 16 48
rect -17 15 -9 18
rect -40 -17 -32 -15
rect -65 -47 -61 -17
rect -35 -47 -32 -17
rect -65 -50 -32 -47
rect -12 -44 -9 15
rect 8 15 16 18
rect 36 44 59 50
rect 8 -44 11 15
rect 36 -15 39 44
rect -12 -50 11 -44
rect 31 -18 39 -15
rect 56 -15 59 44
rect 79 48 112 50
rect 79 18 83 48
rect 109 18 112 48
rect 79 15 87 18
rect 56 -18 64 -15
rect 31 -48 34 -18
rect 60 -48 64 -18
rect 31 -50 64 -48
rect 84 -44 87 15
rect 104 15 112 18
rect 132 44 155 50
rect 104 -44 107 15
rect 132 -15 135 44
rect 84 -50 107 -44
rect 127 -17 135 -15
rect 152 -15 155 44
rect 175 48 208 50
rect 175 18 179 48
rect 205 18 208 48
rect 175 15 183 18
rect 152 -17 160 -15
rect 127 -47 131 -17
rect 157 -47 160 -17
rect 127 -50 160 -47
rect 180 -44 183 15
rect 200 15 208 18
rect 228 44 251 50
rect 200 -44 203 15
rect 228 -15 231 44
rect 180 -50 203 -44
rect 223 -18 231 -15
rect 248 -15 251 44
rect 248 -18 256 -15
rect 223 -48 226 -18
rect 252 -48 256 -18
rect 223 -50 256 -48
rect -39 -69 -10 -66
rect -233 -86 -33 -69
rect -16 -86 223 -69
rect -233 -89 223 -86
<< via1 >>
rect -205 44 -179 48
rect -205 18 -201 44
rect -201 18 -184 44
rect -184 18 -179 44
rect -254 -44 -249 -18
rect -249 -44 -232 -18
rect -232 -44 -228 -18
rect -254 -48 -228 -44
rect -109 44 -83 48
rect -109 18 -105 44
rect -105 18 -88 44
rect -88 18 -83 44
rect -157 -44 -153 -17
rect -153 -44 -136 -17
rect -136 -44 -131 -17
rect -157 -47 -131 -44
rect -14 44 12 48
rect -14 18 -9 44
rect -9 18 8 44
rect 8 18 12 44
rect -61 -44 -57 -17
rect -57 -44 -40 -17
rect -40 -44 -35 -17
rect -61 -47 -35 -44
rect 83 44 109 48
rect 83 18 87 44
rect 87 18 104 44
rect 104 18 109 44
rect 34 -44 39 -18
rect 39 -44 56 -18
rect 56 -44 60 -18
rect 34 -48 60 -44
rect 179 44 205 48
rect 179 18 183 44
rect 183 18 200 44
rect 200 18 205 44
rect 131 -44 135 -17
rect 135 -44 152 -17
rect 152 -44 157 -17
rect 131 -47 157 -44
rect 226 -44 231 -18
rect 231 -44 248 -18
rect 248 -44 252 -18
rect 226 -48 252 -44
<< metal2 >>
rect -257 51 256 94
rect -257 48 133 51
rect -257 18 -205 48
rect -179 18 -109 48
rect -83 18 -14 48
rect 12 18 83 48
rect 109 20 133 48
rect 232 20 256 51
rect 109 18 179 20
rect 205 18 256 20
rect -257 15 256 18
rect -257 -17 256 -15
rect -257 -18 -157 -17
rect -257 -48 -254 -18
rect -228 -21 -157 -18
rect -131 -47 -61 -17
rect -35 -18 131 -17
rect -35 -47 34 -18
rect -143 -48 34 -47
rect 60 -47 131 -18
rect 157 -18 256 -17
rect 157 -47 226 -18
rect 60 -48 226 -47
rect 252 -48 256 -18
rect -257 -52 -242 -48
rect -143 -52 256 -48
rect -257 -94 256 -52
<< via2 >>
rect 133 48 232 51
rect 133 20 179 48
rect 179 20 205 48
rect 205 20 232 48
rect -242 -48 -228 -21
rect -228 -47 -157 -21
rect -157 -47 -143 -21
rect -228 -48 -143 -47
rect -242 -52 -143 -48
<< metal3 >>
rect 124 51 254 59
rect 124 20 133 51
rect 232 20 254 51
rect 124 15 254 20
rect -257 -21 -127 -15
rect -257 -52 -242 -21
rect -143 -52 -127 -21
rect -257 -59 -127 -52
<< properties >>
string FIXED_BBOX -297 -128 297 128
string gencell sky130_fd_pr__nfet_01v8_lvt
string library sky130
string parameters w 1.0 l 0.15 m 1 nf 10 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
