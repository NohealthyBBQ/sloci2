* NGSPICE file created from 3T.ext - technology: sky130A

.subckt sky130_fd_pr__nfet_01v8_lvt_WSE2Y6 a_50_n200# a_n108_n200# a_n50_n288# a_n210_n374#
X0 a_50_n200# a_n50_n288# a_n108_n200# a_n210_n374# sky130_fd_pr__nfet_01v8_lvt ad=5.8e+11p pd=4.58e+06u as=5.8e+11p ps=4.58e+06u w=2e+06u l=500000u
.ends

.subckt sky130_fd_pr__pfet_01v8_LDYTSD a_n50_n297# a_50_n200# a_n108_n200# w_n246_n419#
X0 a_50_n200# a_n50_n297# a_n108_n200# w_n246_n419# sky130_fd_pr__pfet_01v8 ad=5.8e+11p pd=4.58e+06u as=5.8e+11p ps=4.58e+06u w=2e+06u l=500000u
.ends

.subckt 3T Vout rst_b pd_in VDD row_sel VSS
Xsky130_fd_pr__nfet_01v8_lvt_WSE2Y6_0 m1_170_n680# Vout row_sel VSS sky130_fd_pr__nfet_01v8_lvt_WSE2Y6
Xsky130_fd_pr__pfet_01v8_LDYTSD_0 rst_b pd_in VDD VDD sky130_fd_pr__pfet_01v8_LDYTSD
Xsky130_fd_pr__nfet_01v8_lvt_WSE2Y6_1 m1_170_n680# VDD pd_in VSS sky130_fd_pr__nfet_01v8_lvt_WSE2Y6
Xsky130_fd_pr__nfet_01v8_lvt_WSE2Y6_2 m1_170_n680# VDD pd_in VSS sky130_fd_pr__nfet_01v8_lvt_WSE2Y6
.ends

