magic
tech sky130A
magscale 1 2
timestamp 1672261271
<< pwell >>
rect -246 -429 246 429
<< nmoslvt >>
rect -50 -281 50 219
<< ndiff >>
rect -108 207 -50 219
rect -108 -269 -96 207
rect -62 -269 -50 207
rect -108 -281 -50 -269
rect 50 207 108 219
rect 50 -269 62 207
rect 96 -269 108 207
rect 50 -281 108 -269
<< ndiffc >>
rect -96 -269 -62 207
rect 62 -269 96 207
<< psubdiff >>
rect -210 359 210 393
rect -210 297 -176 359
rect 176 297 210 359
rect -210 -359 -176 -297
rect 176 -359 210 -297
rect -210 -393 210 -359
<< psubdiffcont >>
rect -210 -297 -176 297
rect 176 -297 210 297
<< poly >>
rect -50 291 50 307
rect -50 257 -34 291
rect 34 257 50 291
rect -50 219 50 257
rect -50 -307 50 -281
<< polycont >>
rect -34 257 34 291
<< locali >>
rect -210 359 210 393
rect -210 297 -176 359
rect 176 297 210 359
rect -50 257 -34 291
rect 34 257 50 291
rect -96 207 -62 223
rect -96 -285 -62 -269
rect 62 207 96 223
rect 62 -285 96 -269
rect -210 -359 -176 -297
rect 176 -359 210 -297
rect -210 -393 210 -359
<< viali >>
rect -34 257 34 291
rect -96 -269 -62 207
rect 62 -269 96 207
<< metal1 >>
rect -46 291 46 297
rect -46 257 -34 291
rect 34 257 46 291
rect -46 251 46 257
rect -102 207 -56 219
rect -102 -269 -96 207
rect -62 -269 -56 207
rect -102 -281 -56 -269
rect 56 207 102 219
rect 56 -269 62 207
rect 96 -269 102 207
rect 56 -281 102 -269
<< properties >>
string FIXED_BBOX -193 -376 193 376
string gencell sky130_fd_pr__nfet_01v8_lvt
string library sky130
string parameters w 2.5 l 0.5 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 0 gbc 0 tbcov 100 rlcov 100 topc 1 botc 0 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
