magic
tech sky130A
magscale 1 2
timestamp 1672439470
<< psubdiff >>
rect 5870 2040 6008 2078
rect 8908 2040 9204 2078
rect 5870 1934 5904 2040
rect 9170 1924 9204 2040
rect 5870 -386 5904 -198
rect 9170 -354 9204 -208
<< psubdiffcont >>
rect 6008 2040 8908 2078
rect 5870 -198 5904 1934
rect 9170 -208 9204 1924
<< poly >>
rect 6615 1620 6765 1650
rect 6610 1534 6690 1550
rect 6610 1500 6633 1534
rect 6667 1500 6690 1534
rect 6610 1490 6690 1500
rect 6735 1520 6765 1620
rect 6810 1634 6890 1650
rect 6810 1600 6833 1634
rect 6867 1600 6890 1634
rect 7415 1620 7565 1650
rect 6810 1590 6890 1600
rect 7410 1534 7490 1550
rect 6735 1490 6850 1520
rect 7410 1500 7433 1534
rect 7467 1500 7490 1534
rect 7410 1490 7490 1500
rect 7535 1520 7565 1620
rect 7610 1634 7690 1650
rect 7610 1600 7633 1634
rect 7667 1600 7690 1634
rect 8215 1620 8365 1650
rect 7610 1590 7690 1600
rect 8210 1534 8290 1550
rect 7535 1490 7690 1520
rect 8210 1500 8233 1534
rect 8267 1500 8290 1534
rect 8210 1490 8290 1500
rect 8335 1520 8365 1620
rect 8410 1634 8490 1650
rect 8410 1600 8433 1634
rect 8467 1600 8490 1634
rect 8410 1590 8490 1600
rect 8335 1490 8490 1520
rect 6616 1130 6646 1242
rect 6840 1130 6870 1254
rect 7416 1140 7446 1240
rect 7338 1130 7446 1140
rect 7640 1130 7670 1258
rect 8216 1130 8246 1240
rect 8440 1130 8470 1264
rect 6615 1100 6765 1130
rect 6610 1014 6690 1030
rect 6610 980 6633 1014
rect 6667 980 6690 1014
rect 6610 970 6690 980
rect 6735 1000 6765 1100
rect 6810 1114 6890 1130
rect 6810 1080 6833 1114
rect 6867 1080 6890 1114
rect 7338 1124 7565 1130
rect 7338 1090 7361 1124
rect 7395 1100 7565 1124
rect 7395 1090 7418 1100
rect 7338 1080 7418 1090
rect 6810 1070 6890 1080
rect 7410 1014 7490 1030
rect 6735 970 6890 1000
rect 7410 980 7433 1014
rect 7467 980 7490 1014
rect 7410 970 7490 980
rect 7535 1000 7565 1100
rect 7610 1114 7690 1130
rect 7610 1080 7633 1114
rect 7667 1080 7690 1114
rect 8215 1100 8365 1130
rect 7610 1070 7690 1080
rect 8210 1014 8290 1030
rect 7535 970 7690 1000
rect 8210 980 8233 1014
rect 8267 980 8290 1014
rect 8210 970 8290 980
rect 8335 1000 8365 1100
rect 8410 1114 8490 1130
rect 8410 1080 8433 1114
rect 8467 1080 8490 1114
rect 8410 1070 8490 1080
rect 8335 970 8490 1000
rect 6615 680 6765 710
rect 6610 594 6690 610
rect 6610 560 6633 594
rect 6667 560 6690 594
rect 6610 550 6690 560
rect 6735 580 6765 680
rect 6810 694 6890 710
rect 6810 660 6833 694
rect 6867 660 6890 694
rect 7415 680 7565 710
rect 6810 650 6890 660
rect 7410 594 7490 610
rect 6735 550 6890 580
rect 7410 560 7433 594
rect 7467 560 7490 594
rect 7410 550 7490 560
rect 7535 580 7565 680
rect 7610 694 7690 710
rect 7610 660 7633 694
rect 7667 660 7690 694
rect 8215 680 8365 710
rect 7610 650 7690 660
rect 8210 594 8290 610
rect 7535 550 7690 580
rect 8210 560 8233 594
rect 8267 560 8290 594
rect 8210 550 8290 560
rect 8335 580 8365 680
rect 8410 694 8490 710
rect 8410 660 8433 694
rect 8467 660 8490 694
rect 8410 650 8490 660
rect 8335 550 8490 580
rect 6616 190 6646 302
rect 6840 190 6870 314
rect 7416 190 7446 300
rect 7640 190 7670 314
rect 8216 190 8246 300
rect 8440 190 8470 316
rect 6615 160 6765 190
rect 6610 74 6690 90
rect 6610 40 6633 74
rect 6667 40 6690 74
rect 6610 30 6690 40
rect 6735 60 6765 160
rect 6810 174 6890 190
rect 6810 140 6833 174
rect 6867 140 6890 174
rect 7415 160 7565 190
rect 6810 130 6890 140
rect 7410 74 7490 90
rect 6735 30 6890 60
rect 7410 40 7433 74
rect 7467 40 7490 74
rect 7410 30 7490 40
rect 7535 60 7565 160
rect 7610 174 7690 190
rect 7610 140 7633 174
rect 7667 140 7690 174
rect 8215 160 8365 190
rect 7610 130 7690 140
rect 8210 74 8290 90
rect 7535 30 7690 60
rect 8210 40 8233 74
rect 8267 40 8290 74
rect 8210 30 8290 40
rect 8335 60 8365 160
rect 8410 174 8490 190
rect 8410 140 8433 174
rect 8467 140 8490 174
rect 8410 130 8490 140
rect 8335 30 8490 60
<< polycont >>
rect 6633 1500 6667 1534
rect 6833 1600 6867 1634
rect 7433 1500 7467 1534
rect 7633 1600 7667 1634
rect 8233 1500 8267 1534
rect 8433 1600 8467 1634
rect 6633 980 6667 1014
rect 6833 1080 6867 1114
rect 7361 1090 7395 1124
rect 7433 980 7467 1014
rect 7633 1080 7667 1114
rect 8233 980 8267 1014
rect 8433 1080 8467 1114
rect 6633 560 6667 594
rect 6833 660 6867 694
rect 7433 560 7467 594
rect 7633 660 7667 694
rect 8233 560 8267 594
rect 8433 660 8467 694
rect 6633 40 6667 74
rect 6833 140 6867 174
rect 7433 40 7467 74
rect 7633 140 7667 174
rect 8233 40 8267 74
rect 8433 140 8467 174
<< locali >>
rect 7224 2958 7260 3146
rect 7154 2930 7260 2958
rect 7154 2846 7190 2930
rect 7224 2878 7260 2930
rect 7832 3102 7868 3144
rect 7832 3090 7908 3102
rect 7832 3008 7846 3090
rect 7890 3008 7908 3090
rect 7832 2996 7908 3008
rect 7224 2846 7256 2878
rect 7832 2876 7868 2996
rect 7154 2820 7256 2846
rect 7090 2078 7132 2404
rect 7988 2078 8030 2412
rect 5870 2040 6008 2078
rect 8908 2040 9204 2078
rect 5870 1934 5904 2040
rect 9170 1924 9204 2040
rect 6817 1600 6833 1634
rect 6867 1600 6883 1634
rect 7617 1600 7633 1634
rect 7667 1600 7683 1634
rect 8417 1600 8433 1634
rect 8467 1600 8483 1634
rect 6617 1500 6633 1534
rect 6667 1500 6683 1534
rect 7417 1500 7433 1534
rect 7467 1500 7483 1534
rect 8217 1500 8233 1534
rect 8267 1500 8283 1534
rect 6817 1080 6833 1114
rect 6867 1080 6883 1114
rect 7345 1090 7361 1124
rect 7395 1090 7411 1124
rect 7617 1080 7633 1114
rect 7667 1080 7683 1114
rect 8417 1080 8433 1114
rect 8467 1080 8483 1114
rect 6617 980 6633 1014
rect 6667 980 6683 1014
rect 7417 980 7433 1014
rect 7467 980 7483 1014
rect 8217 980 8233 1014
rect 8267 980 8283 1014
rect 6817 660 6833 694
rect 6867 660 6883 694
rect 7617 660 7633 694
rect 7667 660 7683 694
rect 8417 660 8433 694
rect 8467 660 8483 694
rect 6617 560 6633 594
rect 6667 560 6683 594
rect 7417 560 7433 594
rect 7467 560 7483 594
rect 8217 560 8233 594
rect 8267 560 8283 594
rect 6817 140 6833 174
rect 6867 140 6883 174
rect 7617 140 7633 174
rect 7667 140 7683 174
rect 8417 140 8433 174
rect 8467 140 8483 174
rect 6617 40 6633 74
rect 6667 40 6683 74
rect 7417 40 7433 74
rect 7467 40 7483 74
rect 8217 40 8233 74
rect 8267 40 8283 74
rect 5870 -386 5904 -198
rect 7222 -386 7860 -352
rect 9170 -354 9204 -208
rect 7220 -938 7256 -862
rect 7150 -968 7256 -938
rect 7150 -1044 7190 -968
rect 7230 -1006 7256 -968
rect 7826 -950 7862 -862
rect 7826 -982 7912 -950
rect 7230 -1044 7254 -1006
rect 7150 -1074 7254 -1044
rect 7826 -1062 7844 -982
rect 7880 -1062 7912 -982
rect 7826 -1088 7912 -1062
<< viali >>
rect 7190 2846 7224 2930
rect 7846 3008 7890 3090
rect 6833 1600 6867 1634
rect 7633 1600 7667 1634
rect 8433 1600 8467 1634
rect 6633 1500 6667 1534
rect 7433 1500 7467 1534
rect 8233 1500 8267 1534
rect 6833 1080 6867 1114
rect 7361 1090 7395 1124
rect 7633 1080 7667 1114
rect 8433 1080 8467 1114
rect 6633 980 6667 1014
rect 7433 980 7467 1014
rect 8233 980 8267 1014
rect 6833 660 6867 694
rect 7633 660 7667 694
rect 8433 660 8467 694
rect 6633 560 6667 594
rect 7433 560 7467 594
rect 8233 560 8267 594
rect 6833 140 6867 174
rect 7633 140 7667 174
rect 8433 140 8467 174
rect 6633 40 6667 74
rect 7433 40 7467 74
rect 8233 40 8267 74
rect 7190 -1044 7230 -968
rect 7844 -1062 7880 -982
<< metal1 >>
rect 7092 3402 8002 3462
rect 7154 2950 7256 2958
rect 7154 2836 7172 2950
rect 7244 2836 7256 2950
rect 7154 2820 7256 2836
rect 7520 2518 7590 3402
rect 7834 3090 7908 3102
rect 7834 3008 7846 3090
rect 7900 3008 7908 3090
rect 7834 2996 7908 3008
rect 5202 2510 5275 2515
rect 5202 2455 5280 2510
rect 7086 2470 8006 2518
rect 7115 2458 7980 2470
rect 5225 -430 5280 2455
rect 6720 1634 6887 1650
rect 6720 1600 6833 1634
rect 6867 1600 6887 1634
rect 6720 1590 6887 1600
rect 7520 1634 7687 1650
rect 7520 1600 7633 1634
rect 7667 1600 7687 1634
rect 7520 1590 7687 1600
rect 8320 1634 8487 1650
rect 8320 1600 8433 1634
rect 8467 1600 8487 1634
rect 8320 1590 8487 1600
rect 6720 1550 6775 1590
rect 7520 1550 7575 1590
rect 8320 1550 8375 1590
rect 6612 1534 6775 1550
rect 6612 1500 6633 1534
rect 6667 1500 6775 1534
rect 6612 1490 6775 1500
rect 7412 1534 7575 1550
rect 7412 1500 7433 1534
rect 7467 1500 7575 1534
rect 7412 1490 7575 1500
rect 8212 1534 8375 1550
rect 8212 1500 8233 1534
rect 8267 1500 8375 1534
rect 8212 1490 8375 1500
rect 7336 1138 7454 1140
rect 6720 1114 6887 1130
rect 6720 1080 6833 1114
rect 6867 1080 6887 1114
rect 7336 1086 7346 1138
rect 7412 1086 7454 1138
rect 7336 1080 7454 1086
rect 7520 1114 7687 1130
rect 7520 1080 7633 1114
rect 7667 1080 7687 1114
rect 6720 1070 6887 1080
rect 7520 1070 7687 1080
rect 8320 1114 8487 1130
rect 8320 1080 8433 1114
rect 8467 1080 8487 1114
rect 8320 1070 8487 1080
rect 6720 1030 6775 1070
rect 7520 1030 7686 1070
rect 8320 1030 8375 1070
rect 6612 1014 6775 1030
rect 6612 980 6633 1014
rect 6667 980 6775 1014
rect 6612 970 6775 980
rect 7412 1028 7686 1030
rect 7412 1014 7582 1028
rect 7412 980 7433 1014
rect 7467 980 7582 1014
rect 7412 976 7582 980
rect 7678 976 7686 1028
rect 7412 970 7686 976
rect 8212 1014 8375 1030
rect 8212 980 8233 1014
rect 8267 980 8375 1014
rect 8212 970 8375 980
rect 6720 694 6887 710
rect 6720 660 6833 694
rect 6867 660 6887 694
rect 6720 650 6887 660
rect 7520 694 7687 710
rect 7520 660 7633 694
rect 7667 660 7687 694
rect 7520 650 7687 660
rect 8320 694 8487 710
rect 8320 660 8433 694
rect 8467 660 8487 694
rect 8320 650 8487 660
rect 6720 610 6775 650
rect 7520 610 7575 650
rect 8320 610 8375 650
rect 6612 594 6775 610
rect 6612 560 6633 594
rect 6667 560 6775 594
rect 6612 550 6775 560
rect 7412 594 7575 610
rect 7412 560 7433 594
rect 7467 560 7575 594
rect 7412 550 7575 560
rect 8212 594 8375 610
rect 8212 560 8233 594
rect 8267 560 8375 594
rect 8212 550 8375 560
rect 6720 174 6887 190
rect 6720 140 6833 174
rect 6867 140 6887 174
rect 6720 130 6887 140
rect 7520 174 7687 190
rect 7520 140 7633 174
rect 7667 140 7687 174
rect 7520 130 7687 140
rect 8320 174 8487 190
rect 8320 140 8433 174
rect 8467 140 8487 174
rect 8320 130 8487 140
rect 6720 90 6775 130
rect 7520 90 7575 130
rect 8320 90 8375 130
rect 6612 74 6775 90
rect 6612 40 6633 74
rect 6667 40 6775 74
rect 6612 30 6775 40
rect 7412 74 7575 90
rect 7412 40 7433 74
rect 7467 40 7575 74
rect 7412 30 7575 40
rect 8212 74 8375 90
rect 8212 40 8233 74
rect 8267 40 8375 74
rect 8212 30 8375 40
rect 5222 -490 5295 -430
rect 7088 -494 8008 -434
rect 7150 -954 7254 -938
rect 7150 -1054 7174 -954
rect 7236 -1054 7254 -954
rect 7150 -1074 7254 -1054
rect 7510 -1378 7580 -494
rect 7826 -972 7912 -950
rect 7826 -1070 7836 -972
rect 7888 -1070 7912 -972
rect 7826 -1088 7912 -1070
rect 7082 -1438 8012 -1378
rect 7504 -1790 7574 -1438
<< via1 >>
rect 7172 2930 7244 2950
rect 7172 2846 7190 2930
rect 7190 2846 7224 2930
rect 7224 2846 7244 2930
rect 7172 2836 7244 2846
rect 7846 3008 7890 3090
rect 7890 3008 7900 3090
rect 7346 1124 7412 1138
rect 7346 1090 7361 1124
rect 7361 1090 7395 1124
rect 7395 1090 7412 1124
rect 7346 1086 7412 1090
rect 7582 976 7678 1028
rect 7174 -968 7236 -954
rect 7174 -1044 7190 -968
rect 7190 -1044 7230 -968
rect 7230 -1044 7236 -968
rect 7174 -1054 7236 -1044
rect 7836 -982 7888 -972
rect 7836 -1062 7844 -982
rect 7844 -1062 7880 -982
rect 7880 -1062 7888 -982
rect 7836 -1070 7888 -1062
<< metal2 >>
rect 8800 3392 9088 3424
rect 5800 3120 6450 3155
rect 5800 2840 5840 3120
rect 6420 2840 6450 3120
rect 7834 3090 7962 3132
rect 7834 3008 7846 3090
rect 7900 3008 7962 3090
rect 7834 2996 7962 3008
rect 8640 3100 9290 3165
rect 5800 2770 6450 2840
rect 7102 2950 7256 2958
rect 7102 2836 7172 2950
rect 7244 2836 7256 2950
rect 7102 2820 7256 2836
rect 8640 2820 8680 3100
rect 9260 2820 9290 3100
rect 8640 2780 9290 2820
rect 5856 2592 6140 2600
rect 5970 2130 8315 2135
rect 5970 2065 7420 2130
rect 7775 2065 8315 2130
rect 5970 1970 8315 2065
rect 5970 1810 6715 1970
rect 7570 1810 8315 1970
rect 5970 1325 6715 1330
rect 5970 1265 6275 1325
rect 6410 1265 6715 1325
rect 5970 1170 6715 1265
rect 6770 1325 7515 1330
rect 6770 1265 7075 1325
rect 7210 1265 7515 1325
rect 6770 1170 7515 1265
rect 7570 1325 8315 1330
rect 7570 1265 7875 1325
rect 8010 1265 8315 1325
rect 7570 1170 8315 1265
rect 8370 1325 9115 1330
rect 8370 1265 8675 1325
rect 8810 1265 9115 1325
rect 8370 1170 9115 1265
rect 6770 1140 6880 1170
rect 7570 1140 7680 1170
rect 8370 1140 8480 1170
rect 6605 1060 6880 1140
rect 7336 1138 7680 1140
rect 7336 1086 7346 1138
rect 7412 1086 7680 1138
rect 7336 1060 7680 1086
rect 8205 1060 8480 1140
rect 6605 1030 6715 1060
rect 7336 1030 7515 1060
rect 8205 1030 8315 1060
rect 5970 935 6715 1030
rect 5970 875 6270 935
rect 6405 875 6715 935
rect 5970 870 6715 875
rect 6770 935 7515 1030
rect 6770 875 7070 935
rect 7205 875 7515 935
rect 6770 870 7515 875
rect 7570 1028 8315 1030
rect 7570 976 7582 1028
rect 7678 976 8315 1028
rect 7570 935 8315 976
rect 7570 875 7870 935
rect 8005 875 8315 935
rect 7570 870 8315 875
rect 8370 935 9115 1030
rect 8370 875 8670 935
rect 8805 875 9115 935
rect 8370 870 9115 875
rect 5970 385 6715 390
rect 5970 325 6275 385
rect 6410 325 6715 385
rect 5970 230 6715 325
rect 6770 385 7515 390
rect 6770 325 7075 385
rect 7210 325 7515 385
rect 6770 230 7515 325
rect 7570 385 8315 390
rect 7570 325 7875 385
rect 8010 325 8315 385
rect 7570 230 8315 325
rect 8370 385 9115 390
rect 8370 325 8675 385
rect 8810 325 9115 385
rect 8370 230 9115 325
rect 6770 200 6880 230
rect 7570 200 7680 230
rect 8370 200 8480 230
rect 6605 120 6880 200
rect 7405 120 7680 200
rect 8205 120 8480 200
rect 6605 90 6715 120
rect 7405 90 7515 120
rect 8205 90 8315 120
rect 5970 -5 6715 90
rect 5970 -65 6270 -5
rect 6405 -65 6715 -5
rect 5970 -70 6715 -65
rect 6770 -5 7515 90
rect 6770 -65 7070 -5
rect 7205 -65 7515 -5
rect 6770 -70 7515 -65
rect 7570 -5 8315 90
rect 7570 -65 7870 -5
rect 8005 -65 8315 -5
rect 7570 -70 8315 -65
rect 8370 -5 9115 90
rect 8370 -65 8670 -5
rect 8805 -65 9115 -5
rect 8370 -70 9115 -65
rect 5790 -780 6440 -730
rect 5790 -1060 5840 -780
rect 6420 -1060 6440 -780
rect 8625 -780 9275 -735
rect 5790 -1115 6440 -1060
rect 7070 -954 7254 -938
rect 7070 -1054 7174 -954
rect 7236 -1054 7254 -954
rect 7070 -1074 7254 -1054
rect 7826 -972 7972 -950
rect 7826 -1070 7836 -972
rect 7888 -1070 7972 -972
rect 7826 -1088 7972 -1070
rect 8625 -1060 8660 -780
rect 9240 -1060 9275 -780
rect 8625 -1120 9275 -1060
<< via2 >>
rect 5408 3328 6464 3392
rect 8640 3328 9696 3392
rect 5845 3325 6115 3328
rect 5840 2840 6420 3120
rect 8680 2820 9260 3100
rect 5376 2528 6432 2592
rect 8576 2528 9632 2592
rect 8830 2525 9100 2528
rect 7420 2065 7775 2130
rect 7075 1815 7210 1875
rect 8770 1815 8905 1875
rect 6270 1685 6405 1745
rect 7075 1685 7210 1745
rect 7870 1685 8005 1745
rect 8770 1685 8905 1745
rect 6275 1395 6410 1455
rect 7075 1395 7210 1455
rect 7865 1395 8000 1455
rect 8770 1395 8905 1455
rect 6275 1265 6410 1325
rect 7075 1265 7210 1325
rect 7875 1265 8010 1325
rect 8675 1265 8810 1325
rect 6270 875 6405 935
rect 7070 875 7205 935
rect 7870 875 8005 935
rect 8670 875 8805 935
rect 6270 745 6405 805
rect 7075 745 7210 805
rect 7870 745 8005 805
rect 8770 745 8905 805
rect 6275 455 6410 515
rect 7075 455 7210 515
rect 7865 455 8000 515
rect 8770 455 8905 515
rect 6275 325 6410 385
rect 7075 325 7210 385
rect 7875 325 8010 385
rect 8675 325 8810 385
rect 6270 -65 6405 -5
rect 7070 -65 7205 -5
rect 7870 -65 8005 -5
rect 8670 -65 8805 -5
rect 6270 -195 6405 -135
rect 7075 -195 7210 -135
rect 7870 -195 8005 -135
rect 8770 -195 8905 -135
rect 5520 -560 6560 -480
rect 8520 -560 9540 -480
rect 5840 -1060 6420 -780
rect 8660 -1060 9240 -780
rect 5320 -1360 6340 -1280
rect 8500 -1380 9520 -1300
<< metal3 >>
rect 5040 3392 6592 3715
rect 5040 3328 5408 3392
rect 6464 3328 6592 3392
rect 5040 3325 5845 3328
rect 6115 3325 6592 3328
rect 5040 3305 6592 3325
rect 5040 2620 5425 3305
rect 7360 3165 7760 3860
rect 8480 3392 10045 3715
rect 8480 3328 8640 3392
rect 9696 3328 10045 3392
rect 8480 3305 10045 3328
rect 5550 3120 9525 3165
rect 5550 2840 5840 3120
rect 6420 3100 9525 3120
rect 6420 2840 8680 3100
rect 5550 2820 8680 2840
rect 9260 2820 9525 3100
rect 5550 2765 9525 2820
rect 9660 2620 10045 3305
rect 5040 2592 6624 2620
rect 5040 2528 5376 2592
rect 6432 2528 6624 2592
rect 5040 2220 6624 2528
rect 8512 2592 10045 2620
rect 8512 2528 8576 2592
rect 9632 2528 10045 2592
rect 8512 2525 8830 2528
rect 9100 2525 10045 2528
rect 8512 2220 10045 2525
rect 5040 1750 5815 2220
rect 7394 2152 8020 2160
rect 7394 2130 7634 2152
rect 7394 2065 7420 2130
rect 7394 2064 7634 2065
rect 8010 2064 8020 2152
rect 7394 2050 8020 2064
rect 6775 1955 9105 1980
rect 6775 1835 6995 1955
rect 7315 1875 9105 1955
rect 7315 1835 8770 1875
rect 6775 1815 7075 1835
rect 7210 1815 8770 1835
rect 8905 1815 9105 1875
rect 6775 1810 9105 1815
rect 9270 1750 10045 2220
rect 5040 1745 7255 1750
rect 5040 1685 6270 1745
rect 6405 1685 7075 1745
rect 7210 1685 7255 1745
rect 5040 1455 7255 1685
rect 5040 1395 6275 1455
rect 6410 1395 7075 1455
rect 7210 1395 7255 1455
rect 5040 1390 7255 1395
rect 7830 1745 10045 1750
rect 7830 1685 7870 1745
rect 8005 1685 8770 1745
rect 8905 1685 10045 1745
rect 7830 1455 10045 1685
rect 7830 1395 7865 1455
rect 8000 1395 8770 1455
rect 8905 1395 10045 1455
rect 7830 1390 10045 1395
rect 5040 810 5815 1390
rect 6135 1325 6825 1330
rect 6135 1265 6275 1325
rect 6410 1265 6825 1325
rect 6135 1160 6825 1265
rect 6935 1325 7625 1330
rect 6935 1265 7075 1325
rect 7210 1265 7625 1325
rect 6935 1160 7625 1265
rect 7735 1325 8420 1330
rect 7735 1265 7875 1325
rect 8010 1265 8420 1325
rect 7735 1160 8420 1265
rect 8535 1325 9115 1330
rect 8535 1265 8675 1325
rect 8810 1265 9115 1325
rect 8535 1160 9115 1265
rect 6660 1040 6825 1160
rect 7460 1040 7625 1160
rect 8255 1040 8420 1160
rect 5970 935 6550 1040
rect 5970 875 6270 935
rect 6405 875 6550 935
rect 5970 870 6550 875
rect 6660 1020 7350 1040
rect 6660 900 6985 1020
rect 7305 900 7350 1020
rect 6660 875 7070 900
rect 7205 875 7350 900
rect 6660 870 7350 875
rect 7460 1010 8150 1040
rect 7460 890 7655 1010
rect 7975 935 8150 1010
rect 7460 875 7870 890
rect 8005 875 8150 935
rect 7460 870 8150 875
rect 8255 935 8950 1040
rect 8255 875 8670 935
rect 8805 875 8950 935
rect 8255 870 8950 875
rect 9270 810 10045 1390
rect 5040 805 7255 810
rect 5040 745 6270 805
rect 6405 745 7075 805
rect 7210 745 7255 805
rect 5040 515 7255 745
rect 5040 455 6275 515
rect 6410 455 7075 515
rect 7210 455 7255 515
rect 5040 450 7255 455
rect 7830 805 10045 810
rect 7830 745 7870 805
rect 8005 745 8770 805
rect 8905 745 10045 805
rect 7830 515 10045 745
rect 7830 455 7865 515
rect 8000 455 8770 515
rect 8905 455 10045 515
rect 7830 450 10045 455
rect 5040 -130 5815 450
rect 6135 385 6820 390
rect 6135 325 6275 385
rect 6410 325 6820 385
rect 6135 220 6820 325
rect 6935 385 7620 390
rect 6935 325 7075 385
rect 7210 325 7620 385
rect 6935 220 7620 325
rect 7735 385 8425 390
rect 7735 325 7875 385
rect 8010 325 8425 385
rect 7735 220 8425 325
rect 8535 385 9115 390
rect 8535 325 8675 385
rect 8810 325 9115 385
rect 8535 220 9115 325
rect 6655 100 6820 220
rect 7455 100 7620 220
rect 8260 100 8425 220
rect 5970 -5 6550 100
rect 5970 -65 6270 -5
rect 6405 -65 6550 -5
rect 5970 -70 6550 -65
rect 6655 80 7350 100
rect 6655 -40 6990 80
rect 7310 -40 7350 80
rect 6655 -65 7070 -40
rect 7205 -65 7350 -40
rect 6655 -70 7350 -65
rect 7455 75 8150 100
rect 7455 -45 7660 75
rect 7980 -5 8150 75
rect 7455 -65 7870 -45
rect 8005 -65 8150 -5
rect 7455 -70 8150 -65
rect 8260 -5 8950 100
rect 8260 -65 8670 -5
rect 8805 -65 8950 -5
rect 8260 -70 8950 -65
rect 9270 -130 10045 450
rect 5040 -135 10045 -130
rect 5040 -195 6270 -135
rect 6405 -195 7075 -135
rect 7210 -195 7870 -135
rect 8005 -195 8770 -135
rect 8905 -195 10045 -135
rect 5040 -480 10045 -195
rect 5040 -560 5520 -480
rect 6560 -560 8520 -480
rect 9540 -560 10045 -480
rect 5040 -575 10045 -560
rect 5040 -1275 5425 -575
rect 5550 -780 9525 -735
rect 5550 -1060 5840 -780
rect 6420 -1060 8660 -780
rect 9240 -1060 9525 -780
rect 5550 -1135 9525 -1060
rect 5040 -1280 6620 -1275
rect 5040 -1360 5320 -1280
rect 6340 -1360 6620 -1280
rect 5040 -1675 6620 -1360
rect 7260 -1780 7780 -1135
rect 9660 -1275 10045 -575
rect 8380 -1300 10045 -1275
rect 8380 -1380 8500 -1300
rect 9520 -1380 10045 -1300
rect 8380 -1675 10045 -1380
<< via3 >>
rect 7634 2130 8010 2152
rect 7634 2065 7775 2130
rect 7775 2065 8010 2130
rect 7634 2064 8010 2065
rect 6995 1875 7315 1955
rect 6995 1835 7075 1875
rect 7075 1835 7210 1875
rect 7210 1835 7315 1875
rect 6985 935 7305 1020
rect 6985 900 7070 935
rect 7070 900 7205 935
rect 7205 900 7305 935
rect 7655 935 7975 1010
rect 7655 890 7870 935
rect 7870 890 7975 935
rect 6990 -5 7310 80
rect 6990 -40 7070 -5
rect 7070 -40 7205 -5
rect 7205 -40 7310 -5
rect 7660 -5 7980 75
rect 7660 -45 7870 -5
rect 7870 -45 7980 -5
<< metal4 >>
rect 7620 2152 8020 2160
rect 7620 2064 7634 2152
rect 8010 2064 8020 2152
rect 6945 1955 7350 1985
rect 6945 1835 6995 1955
rect 7315 1835 7350 1955
rect 6945 1740 7350 1835
rect 3440 1700 7350 1740
rect 3440 1460 3480 1700
rect 3720 1460 7350 1700
rect 3440 1420 7350 1460
rect 6945 1020 7350 1420
rect 6945 900 6985 1020
rect 7305 900 7350 1020
rect 6945 80 7350 900
rect 6945 -40 6990 80
rect 7310 -40 7350 80
rect 6945 -70 7350 -40
rect 7620 1740 8020 2064
rect 7620 1700 11540 1740
rect 7620 1460 11230 1700
rect 11470 1460 11540 1700
rect 7620 1420 11540 1460
rect 7620 1010 8020 1420
rect 7620 890 7655 1010
rect 7975 890 8020 1010
rect 7620 75 8020 890
rect 7620 -45 7660 75
rect 7980 -45 8020 75
rect 7620 -70 8020 -45
<< via4 >>
rect 3480 1460 3720 1700
rect 11230 1460 11470 1700
<< metal5 >>
rect 1520 3340 6320 3660
rect 1520 -180 1840 3340
rect 2160 2700 5680 3020
rect 2160 460 2480 2700
rect 2800 2060 5040 2380
rect 2800 1100 3120 2060
rect 3440 1700 4400 1740
rect 3440 1460 3480 1700
rect 3720 1460 4400 1700
rect 3440 1420 4400 1460
rect 4080 1100 4400 1420
rect 2800 780 4400 1100
rect 4720 460 5040 2060
rect 2160 140 5040 460
rect 5360 -180 5680 2700
rect 1520 -500 5680 -180
rect 6000 -820 6320 3340
rect 9270 3340 14070 3660
rect 9270 -180 9590 3340
rect 9910 2700 13430 3020
rect 9910 460 10230 2700
rect 10550 2060 12790 2380
rect 10550 1100 10870 2060
rect 11190 1700 12150 1740
rect 11190 1460 11230 1700
rect 11470 1460 12150 1700
rect 11190 1420 12150 1460
rect 11830 1100 12150 1420
rect 10550 780 12150 1100
rect 12470 460 12790 2060
rect 9910 140 12790 460
rect 13110 -180 13430 2700
rect 9270 -500 13430 -180
rect 13750 -820 14070 3340
rect 1520 -832 6320 -820
rect 1504 -1140 6320 -832
rect 9270 -1140 14070 -820
rect 1504 -1632 1856 -1140
rect 9280 -1632 9632 -1140
use sky130_fd_pr__nfet_01v8_lvt_WKNS5B  XM1
timestamp 1671055274
transform 1 0 7123 0 1 1770
box -480 -300 526 320
use sky130_fd_pr__nfet_01v8_lvt_WKNS5B  XM2
timestamp 1671055274
transform 1 0 7920 0 1 1350
box -480 -300 526 320
use sky130_fd_pr__nfet_01v8_lvt_WKNS5B  XM3
timestamp 1671055274
transform 1 0 7120 0 1 830
box -480 -300 526 320
use sky130_fd_pr__nfet_01v8_lvt_WKNS5B  XM4
timestamp 1671055274
transform 1 0 7920 0 1 410
box -480 -300 526 320
use sky130_fd_pr__nfet_01v8_lvt_WKNS5B  XM5
timestamp 1671055274
transform 1 0 7120 0 1 -110
box -480 -300 526 320
use sky130_fd_pr__nfet_01v8_lvt_WKNS5B  XM6
timestamp 1671055274
transform 1 0 8720 0 1 1770
box -480 -300 526 320
use sky130_fd_pr__nfet_01v8_lvt_WKNS5B  XM7
timestamp 1671055274
transform 1 0 6320 0 1 1350
box -480 -300 526 320
use sky130_fd_pr__nfet_01v8_lvt_WKNS5B  XM8
timestamp 1671055274
transform 1 0 8720 0 1 830
box -480 -300 526 320
use sky130_fd_pr__nfet_01v8_lvt_WKNS5B  XM9
timestamp 1671055274
transform 1 0 8720 0 1 410
box -480 -300 526 320
use sky130_fd_pr__nfet_01v8_lvt_WKNS5B  XM10
timestamp 1671055274
transform 1 0 6320 0 1 -110
box -480 -300 526 320
use sky130_fd_pr__nfet_01v8_lvt_WKNS5B  XM11
timestamp 1671055274
transform 1 0 7920 0 1 1770
box -480 -300 526 320
use sky130_fd_pr__nfet_01v8_lvt_WKNS5B  XM12
timestamp 1671055274
transform 1 0 7120 0 1 1350
box -480 -300 526 320
use sky130_fd_pr__nfet_01v8_lvt_WKNS5B  XM13
timestamp 1671055274
transform 1 0 7920 0 1 830
box -480 -300 526 320
use sky130_fd_pr__nfet_01v8_lvt_WKNS5B  XM14
timestamp 1671055274
transform 1 0 7120 0 1 410
box -480 -300 526 320
use sky130_fd_pr__nfet_01v8_lvt_WKNS5B  XM15
timestamp 1671055274
transform 1 0 7920 0 1 -110
box -480 -300 526 320
use sky130_fd_pr__nfet_01v8_lvt_WKNS5B  XM16
timestamp 1671055274
transform 1 0 6320 0 1 1770
box -480 -300 526 320
use sky130_fd_pr__nfet_01v8_lvt_WKNS5B  XM17
timestamp 1671055274
transform 1 0 8720 0 1 1350
box -480 -300 526 320
use sky130_fd_pr__nfet_01v8_lvt_WKNS5B  XM18
timestamp 1671055274
transform 1 0 6320 0 1 830
box -480 -300 526 320
use sky130_fd_pr__nfet_01v8_lvt_WKNS5B  XM19
timestamp 1671055274
transform -1 0 6366 0 1 410
box -480 -300 526 320
use sky130_fd_pr__nfet_01v8_lvt_YTLFGX#0  XM21
timestamp 1671827388
transform 1 0 6168 0 1 2650
box -1128 -310 1126 310
use sky130_fd_pr__nfet_01v8_lvt_YTLFGX#0  XM22
timestamp 1671827388
transform -1 0 8922 0 1 2650
box -1128 -310 1126 310
use sky130_fd_pr__nfet_01v8_lvt_YTLFGX#0  XM23
timestamp 1671827388
transform 1 0 6166 0 -1 -626
box -1128 -310 1126 310
use sky130_fd_pr__nfet_01v8_lvt_YTLFGX#0  XM24
timestamp 1671827388
transform -1 0 8916 0 -1 -626
box -1128 -310 1126 310
use sky130_fd_pr__nfet_01v8_lvt_YTLFGX#0  XM25
timestamp 1671827388
transform 1 0 6168 0 -1 3270
box -1128 -310 1126 310
use sky130_fd_pr__nfet_01v8_lvt_YTLFGX#0  XM26
timestamp 1671827388
transform -1 0 8922 0 -1 3270
box -1128 -310 1126 310
use sky130_fd_pr__nfet_01v8_lvt_YTLFGX#0  XM27
timestamp 1671827388
transform 1 0 6166 0 1 -1246
box -1128 -310 1126 310
use sky130_fd_pr__nfet_01v8_lvt_YTLFGX#0  XM28
timestamp 1671827388
transform -1 0 8916 0 1 -1246
box -1128 -310 1126 310
use sky130_fd_pr__nfet_01v8_lvt_WKNS5B  sky130_fd_pr__nfet_01v8_lvt_WKNS5B_1
timestamp 1671055274
transform 1 0 8720 0 1 -110
box -480 -300 526 320
<< labels >>
flabel metal4 7620 1420 11230 1740 0 FreeSans 1600 0 0 0 cap2
flabel metal4 3720 1420 7350 1740 0 FreeSans 1600 0 0 0 cap1
flabel metal3 7360 3160 7760 3860 0 FreeSans 1600 0 0 0 VSS
flabel metal3 7260 -1780 7780 -1080 0 FreeSans 1600 0 0 0 VSS
<< end >>
