magic
tech sky130A
magscale 1 2
timestamp 1662090071
<< nmoslvt >>
rect -487 -419 -287 481
rect -229 -419 -29 481
rect 29 -419 229 481
rect 287 -419 487 481
<< ndiff >>
rect -545 469 -487 481
rect -545 -407 -533 469
rect -499 -407 -487 469
rect -545 -419 -487 -407
rect -287 469 -229 481
rect -287 -407 -275 469
rect -241 -407 -229 469
rect -287 -419 -229 -407
rect -29 469 29 481
rect -29 -407 -17 469
rect 17 -407 29 469
rect -29 -419 29 -407
rect 229 469 287 481
rect 229 -407 241 469
rect 275 -407 287 469
rect 229 -419 287 -407
rect 487 469 545 481
rect 487 -407 499 469
rect 533 -407 545 469
rect 487 -419 545 -407
<< ndiffc >>
rect -533 -407 -499 469
rect -275 -407 -241 469
rect -17 -407 17 469
rect 241 -407 275 469
rect 499 -407 533 469
<< poly >>
rect -487 481 -287 507
rect -229 481 -29 507
rect 29 481 229 507
rect 287 481 487 507
rect -487 -457 -287 -419
rect -487 -491 -471 -457
rect -303 -491 -287 -457
rect -487 -507 -287 -491
rect -229 -457 -29 -419
rect -229 -491 -213 -457
rect -45 -491 -29 -457
rect -229 -507 -29 -491
rect 29 -457 229 -419
rect 29 -491 45 -457
rect 213 -491 229 -457
rect 29 -507 229 -491
rect 287 -457 487 -419
rect 287 -491 303 -457
rect 471 -491 487 -457
rect 287 -507 487 -491
<< polycont >>
rect -471 -491 -303 -457
rect -213 -491 -45 -457
rect 45 -491 213 -457
rect 303 -491 471 -457
<< locali >>
rect -533 469 -499 485
rect -533 -423 -499 -407
rect -275 469 -241 485
rect -275 -423 -241 -407
rect -17 469 17 485
rect -17 -423 17 -407
rect 241 469 275 485
rect 241 -423 275 -407
rect 499 469 533 485
rect 499 -423 533 -407
rect -487 -491 -471 -457
rect -303 -491 -287 -457
rect -229 -491 -213 -457
rect -45 -491 -29 -457
rect 29 -491 45 -457
rect 213 -491 229 -457
rect 287 -491 303 -457
rect 471 -491 487 -457
<< viali >>
rect -533 -407 -499 469
rect -275 -407 -241 469
rect -17 -407 17 469
rect 241 -407 275 469
rect 499 -407 533 469
rect -471 -491 -303 -457
rect -213 -491 -45 -457
rect 45 -491 213 -457
rect 303 -491 471 -457
<< metal1 >>
rect -539 469 -493 481
rect -539 -407 -533 469
rect -499 -407 -493 469
rect -539 -419 -493 -407
rect -281 469 -235 481
rect -281 -407 -275 469
rect -241 -407 -235 469
rect -281 -419 -235 -407
rect -23 469 23 481
rect -23 -407 -17 469
rect 17 -407 23 469
rect -23 -419 23 -407
rect 235 469 281 481
rect 235 -407 241 469
rect 275 -407 281 469
rect 235 -419 281 -407
rect 493 469 539 481
rect 493 -407 499 469
rect 533 -407 539 469
rect 493 -419 539 -407
rect -483 -457 -291 -451
rect -483 -491 -471 -457
rect -303 -491 -291 -457
rect -483 -497 -291 -491
rect -225 -457 -33 -451
rect -225 -491 -213 -457
rect -45 -491 -33 -457
rect -225 -497 -33 -491
rect 33 -457 225 -451
rect 33 -491 45 -457
rect 213 -491 225 -457
rect 33 -497 225 -491
rect 291 -457 483 -451
rect 291 -491 303 -457
rect 471 -491 483 -457
rect 291 -497 483 -491
<< properties >>
string gencell sky130_fd_pr__nfet_01v8_lvt
string library sky130
string parameters w 4.5 l 1 m 1 nf 4 diffcov 100 polycov 100 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 0 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 0 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
