magic
tech sky130A
magscale 1 2
timestamp 1671745787
<< error_p >>
rect -461 799 -403 805
rect -269 799 -211 805
rect -77 799 -19 805
rect 115 799 173 805
rect 307 799 365 805
rect -461 765 -449 799
rect -269 765 -257 799
rect -77 765 -65 799
rect 115 765 127 799
rect 307 765 319 799
rect -461 759 -403 765
rect -269 759 -211 765
rect -77 759 -19 765
rect 115 759 173 765
rect 307 759 365 765
rect -365 489 -307 495
rect -173 489 -115 495
rect 19 489 77 495
rect 211 489 269 495
rect 403 489 461 495
rect -365 455 -353 489
rect -173 455 -161 489
rect 19 455 31 489
rect 211 455 223 489
rect 403 455 415 489
rect -365 449 -307 455
rect -173 449 -115 455
rect 19 449 77 455
rect 211 449 269 455
rect 403 449 461 455
rect -365 381 -307 387
rect -173 381 -115 387
rect 19 381 77 387
rect 211 381 269 387
rect 403 381 461 387
rect -365 347 -353 381
rect -173 347 -161 381
rect 19 347 31 381
rect 211 347 223 381
rect 403 347 415 381
rect -365 341 -307 347
rect -173 341 -115 347
rect 19 341 77 347
rect 211 341 269 347
rect 403 341 461 347
rect -461 71 -403 77
rect -269 71 -211 77
rect -77 71 -19 77
rect 115 71 173 77
rect 307 71 365 77
rect -461 37 -449 71
rect -269 37 -257 71
rect -77 37 -65 71
rect 115 37 127 71
rect 307 37 319 71
rect -461 31 -403 37
rect -269 31 -211 37
rect -77 31 -19 37
rect 115 31 173 37
rect 307 31 365 37
rect -461 -37 -403 -31
rect -269 -37 -211 -31
rect -77 -37 -19 -31
rect 115 -37 173 -31
rect 307 -37 365 -31
rect -461 -71 -449 -37
rect -269 -71 -257 -37
rect -77 -71 -65 -37
rect 115 -71 127 -37
rect 307 -71 319 -37
rect -461 -77 -403 -71
rect -269 -77 -211 -71
rect -77 -77 -19 -71
rect 115 -77 173 -71
rect 307 -77 365 -71
rect -365 -347 -307 -341
rect -173 -347 -115 -341
rect 19 -347 77 -341
rect 211 -347 269 -341
rect 403 -347 461 -341
rect -365 -381 -353 -347
rect -173 -381 -161 -347
rect 19 -381 31 -347
rect 211 -381 223 -347
rect 403 -381 415 -347
rect -365 -387 -307 -381
rect -173 -387 -115 -381
rect 19 -387 77 -381
rect 211 -387 269 -381
rect 403 -387 461 -381
rect -365 -455 -307 -449
rect -173 -455 -115 -449
rect 19 -455 77 -449
rect 211 -455 269 -449
rect 403 -455 461 -449
rect -365 -489 -353 -455
rect -173 -489 -161 -455
rect 19 -489 31 -455
rect 211 -489 223 -455
rect 403 -489 415 -455
rect -365 -495 -307 -489
rect -173 -495 -115 -489
rect 19 -495 77 -489
rect 211 -495 269 -489
rect 403 -495 461 -489
rect -461 -765 -403 -759
rect -269 -765 -211 -759
rect -77 -765 -19 -759
rect 115 -765 173 -759
rect 307 -765 365 -759
rect -461 -799 -449 -765
rect -269 -799 -257 -765
rect -77 -799 -65 -765
rect 115 -799 127 -765
rect 307 -799 319 -765
rect -461 -805 -403 -799
rect -269 -805 -211 -799
rect -77 -805 -19 -799
rect 115 -805 173 -799
rect 307 -805 365 -799
<< pwell >>
rect -647 -937 647 937
<< nmoslvt >>
rect -447 527 -417 727
rect -351 527 -321 727
rect -255 527 -225 727
rect -159 527 -129 727
rect -63 527 -33 727
rect 33 527 63 727
rect 129 527 159 727
rect 225 527 255 727
rect 321 527 351 727
rect 417 527 447 727
rect -447 109 -417 309
rect -351 109 -321 309
rect -255 109 -225 309
rect -159 109 -129 309
rect -63 109 -33 309
rect 33 109 63 309
rect 129 109 159 309
rect 225 109 255 309
rect 321 109 351 309
rect 417 109 447 309
rect -447 -309 -417 -109
rect -351 -309 -321 -109
rect -255 -309 -225 -109
rect -159 -309 -129 -109
rect -63 -309 -33 -109
rect 33 -309 63 -109
rect 129 -309 159 -109
rect 225 -309 255 -109
rect 321 -309 351 -109
rect 417 -309 447 -109
rect -447 -727 -417 -527
rect -351 -727 -321 -527
rect -255 -727 -225 -527
rect -159 -727 -129 -527
rect -63 -727 -33 -527
rect 33 -727 63 -527
rect 129 -727 159 -527
rect 225 -727 255 -527
rect 321 -727 351 -527
rect 417 -727 447 -527
<< ndiff >>
rect -509 715 -447 727
rect -509 539 -497 715
rect -463 539 -447 715
rect -509 527 -447 539
rect -417 715 -351 727
rect -417 539 -401 715
rect -367 539 -351 715
rect -417 527 -351 539
rect -321 715 -255 727
rect -321 539 -305 715
rect -271 539 -255 715
rect -321 527 -255 539
rect -225 715 -159 727
rect -225 539 -209 715
rect -175 539 -159 715
rect -225 527 -159 539
rect -129 715 -63 727
rect -129 539 -113 715
rect -79 539 -63 715
rect -129 527 -63 539
rect -33 715 33 727
rect -33 539 -17 715
rect 17 539 33 715
rect -33 527 33 539
rect 63 715 129 727
rect 63 539 79 715
rect 113 539 129 715
rect 63 527 129 539
rect 159 715 225 727
rect 159 539 175 715
rect 209 539 225 715
rect 159 527 225 539
rect 255 715 321 727
rect 255 539 271 715
rect 305 539 321 715
rect 255 527 321 539
rect 351 715 417 727
rect 351 539 367 715
rect 401 539 417 715
rect 351 527 417 539
rect 447 715 509 727
rect 447 539 463 715
rect 497 539 509 715
rect 447 527 509 539
rect -509 297 -447 309
rect -509 121 -497 297
rect -463 121 -447 297
rect -509 109 -447 121
rect -417 297 -351 309
rect -417 121 -401 297
rect -367 121 -351 297
rect -417 109 -351 121
rect -321 297 -255 309
rect -321 121 -305 297
rect -271 121 -255 297
rect -321 109 -255 121
rect -225 297 -159 309
rect -225 121 -209 297
rect -175 121 -159 297
rect -225 109 -159 121
rect -129 297 -63 309
rect -129 121 -113 297
rect -79 121 -63 297
rect -129 109 -63 121
rect -33 297 33 309
rect -33 121 -17 297
rect 17 121 33 297
rect -33 109 33 121
rect 63 297 129 309
rect 63 121 79 297
rect 113 121 129 297
rect 63 109 129 121
rect 159 297 225 309
rect 159 121 175 297
rect 209 121 225 297
rect 159 109 225 121
rect 255 297 321 309
rect 255 121 271 297
rect 305 121 321 297
rect 255 109 321 121
rect 351 297 417 309
rect 351 121 367 297
rect 401 121 417 297
rect 351 109 417 121
rect 447 297 509 309
rect 447 121 463 297
rect 497 121 509 297
rect 447 109 509 121
rect -509 -121 -447 -109
rect -509 -297 -497 -121
rect -463 -297 -447 -121
rect -509 -309 -447 -297
rect -417 -121 -351 -109
rect -417 -297 -401 -121
rect -367 -297 -351 -121
rect -417 -309 -351 -297
rect -321 -121 -255 -109
rect -321 -297 -305 -121
rect -271 -297 -255 -121
rect -321 -309 -255 -297
rect -225 -121 -159 -109
rect -225 -297 -209 -121
rect -175 -297 -159 -121
rect -225 -309 -159 -297
rect -129 -121 -63 -109
rect -129 -297 -113 -121
rect -79 -297 -63 -121
rect -129 -309 -63 -297
rect -33 -121 33 -109
rect -33 -297 -17 -121
rect 17 -297 33 -121
rect -33 -309 33 -297
rect 63 -121 129 -109
rect 63 -297 79 -121
rect 113 -297 129 -121
rect 63 -309 129 -297
rect 159 -121 225 -109
rect 159 -297 175 -121
rect 209 -297 225 -121
rect 159 -309 225 -297
rect 255 -121 321 -109
rect 255 -297 271 -121
rect 305 -297 321 -121
rect 255 -309 321 -297
rect 351 -121 417 -109
rect 351 -297 367 -121
rect 401 -297 417 -121
rect 351 -309 417 -297
rect 447 -121 509 -109
rect 447 -297 463 -121
rect 497 -297 509 -121
rect 447 -309 509 -297
rect -509 -539 -447 -527
rect -509 -715 -497 -539
rect -463 -715 -447 -539
rect -509 -727 -447 -715
rect -417 -539 -351 -527
rect -417 -715 -401 -539
rect -367 -715 -351 -539
rect -417 -727 -351 -715
rect -321 -539 -255 -527
rect -321 -715 -305 -539
rect -271 -715 -255 -539
rect -321 -727 -255 -715
rect -225 -539 -159 -527
rect -225 -715 -209 -539
rect -175 -715 -159 -539
rect -225 -727 -159 -715
rect -129 -539 -63 -527
rect -129 -715 -113 -539
rect -79 -715 -63 -539
rect -129 -727 -63 -715
rect -33 -539 33 -527
rect -33 -715 -17 -539
rect 17 -715 33 -539
rect -33 -727 33 -715
rect 63 -539 129 -527
rect 63 -715 79 -539
rect 113 -715 129 -539
rect 63 -727 129 -715
rect 159 -539 225 -527
rect 159 -715 175 -539
rect 209 -715 225 -539
rect 159 -727 225 -715
rect 255 -539 321 -527
rect 255 -715 271 -539
rect 305 -715 321 -539
rect 255 -727 321 -715
rect 351 -539 417 -527
rect 351 -715 367 -539
rect 401 -715 417 -539
rect 351 -727 417 -715
rect 447 -539 509 -527
rect 447 -715 463 -539
rect 497 -715 509 -539
rect 447 -727 509 -715
<< ndiffc >>
rect -497 539 -463 715
rect -401 539 -367 715
rect -305 539 -271 715
rect -209 539 -175 715
rect -113 539 -79 715
rect -17 539 17 715
rect 79 539 113 715
rect 175 539 209 715
rect 271 539 305 715
rect 367 539 401 715
rect 463 539 497 715
rect -497 121 -463 297
rect -401 121 -367 297
rect -305 121 -271 297
rect -209 121 -175 297
rect -113 121 -79 297
rect -17 121 17 297
rect 79 121 113 297
rect 175 121 209 297
rect 271 121 305 297
rect 367 121 401 297
rect 463 121 497 297
rect -497 -297 -463 -121
rect -401 -297 -367 -121
rect -305 -297 -271 -121
rect -209 -297 -175 -121
rect -113 -297 -79 -121
rect -17 -297 17 -121
rect 79 -297 113 -121
rect 175 -297 209 -121
rect 271 -297 305 -121
rect 367 -297 401 -121
rect 463 -297 497 -121
rect -497 -715 -463 -539
rect -401 -715 -367 -539
rect -305 -715 -271 -539
rect -209 -715 -175 -539
rect -113 -715 -79 -539
rect -17 -715 17 -539
rect 79 -715 113 -539
rect 175 -715 209 -539
rect 271 -715 305 -539
rect 367 -715 401 -539
rect 463 -715 497 -539
<< psubdiff >>
rect -611 867 -515 901
rect 515 867 611 901
rect -611 805 -577 867
rect 577 805 611 867
rect -611 -867 -577 -805
rect 577 -867 611 -805
rect -611 -901 -515 -867
rect 515 -901 611 -867
<< psubdiffcont >>
rect -515 867 515 901
rect -611 -805 -577 805
rect 577 -805 611 805
rect -515 -901 515 -867
<< poly >>
rect -465 799 -399 815
rect -465 765 -449 799
rect -415 765 -399 799
rect -465 749 -399 765
rect -273 799 -207 815
rect -273 765 -257 799
rect -223 765 -207 799
rect -447 727 -417 749
rect -351 727 -321 753
rect -273 749 -207 765
rect -81 799 -15 815
rect -81 765 -65 799
rect -31 765 -15 799
rect -255 727 -225 749
rect -159 727 -129 753
rect -81 749 -15 765
rect 111 799 177 815
rect 111 765 127 799
rect 161 765 177 799
rect -63 727 -33 749
rect 33 727 63 753
rect 111 749 177 765
rect 303 799 369 815
rect 303 765 319 799
rect 353 765 369 799
rect 129 727 159 749
rect 225 727 255 753
rect 303 749 369 765
rect 321 727 351 749
rect 417 727 447 753
rect -447 501 -417 527
rect -351 505 -321 527
rect -369 489 -303 505
rect -255 501 -225 527
rect -159 505 -129 527
rect -369 455 -353 489
rect -319 455 -303 489
rect -369 439 -303 455
rect -177 489 -111 505
rect -63 501 -33 527
rect 33 505 63 527
rect -177 455 -161 489
rect -127 455 -111 489
rect -177 439 -111 455
rect 15 489 81 505
rect 129 501 159 527
rect 225 505 255 527
rect 15 455 31 489
rect 65 455 81 489
rect 15 439 81 455
rect 207 489 273 505
rect 321 501 351 527
rect 417 505 447 527
rect 207 455 223 489
rect 257 455 273 489
rect 207 439 273 455
rect 399 489 465 505
rect 399 455 415 489
rect 449 455 465 489
rect 399 439 465 455
rect -369 381 -303 397
rect -369 347 -353 381
rect -319 347 -303 381
rect -447 309 -417 335
rect -369 331 -303 347
rect -177 381 -111 397
rect -177 347 -161 381
rect -127 347 -111 381
rect -351 309 -321 331
rect -255 309 -225 335
rect -177 331 -111 347
rect 15 381 81 397
rect 15 347 31 381
rect 65 347 81 381
rect -159 309 -129 331
rect -63 309 -33 335
rect 15 331 81 347
rect 207 381 273 397
rect 207 347 223 381
rect 257 347 273 381
rect 33 309 63 331
rect 129 309 159 335
rect 207 331 273 347
rect 399 381 465 397
rect 399 347 415 381
rect 449 347 465 381
rect 225 309 255 331
rect 321 309 351 335
rect 399 331 465 347
rect 417 309 447 331
rect -447 87 -417 109
rect -465 71 -399 87
rect -351 83 -321 109
rect -255 87 -225 109
rect -465 37 -449 71
rect -415 37 -399 71
rect -465 21 -399 37
rect -273 71 -207 87
rect -159 83 -129 109
rect -63 87 -33 109
rect -273 37 -257 71
rect -223 37 -207 71
rect -273 21 -207 37
rect -81 71 -15 87
rect 33 83 63 109
rect 129 87 159 109
rect -81 37 -65 71
rect -31 37 -15 71
rect -81 21 -15 37
rect 111 71 177 87
rect 225 83 255 109
rect 321 87 351 109
rect 111 37 127 71
rect 161 37 177 71
rect 111 21 177 37
rect 303 71 369 87
rect 417 83 447 109
rect 303 37 319 71
rect 353 37 369 71
rect 303 21 369 37
rect -465 -37 -399 -21
rect -465 -71 -449 -37
rect -415 -71 -399 -37
rect -465 -87 -399 -71
rect -273 -37 -207 -21
rect -273 -71 -257 -37
rect -223 -71 -207 -37
rect -447 -109 -417 -87
rect -351 -109 -321 -83
rect -273 -87 -207 -71
rect -81 -37 -15 -21
rect -81 -71 -65 -37
rect -31 -71 -15 -37
rect -255 -109 -225 -87
rect -159 -109 -129 -83
rect -81 -87 -15 -71
rect 111 -37 177 -21
rect 111 -71 127 -37
rect 161 -71 177 -37
rect -63 -109 -33 -87
rect 33 -109 63 -83
rect 111 -87 177 -71
rect 303 -37 369 -21
rect 303 -71 319 -37
rect 353 -71 369 -37
rect 129 -109 159 -87
rect 225 -109 255 -83
rect 303 -87 369 -71
rect 321 -109 351 -87
rect 417 -109 447 -83
rect -447 -335 -417 -309
rect -351 -331 -321 -309
rect -369 -347 -303 -331
rect -255 -335 -225 -309
rect -159 -331 -129 -309
rect -369 -381 -353 -347
rect -319 -381 -303 -347
rect -369 -397 -303 -381
rect -177 -347 -111 -331
rect -63 -335 -33 -309
rect 33 -331 63 -309
rect -177 -381 -161 -347
rect -127 -381 -111 -347
rect -177 -397 -111 -381
rect 15 -347 81 -331
rect 129 -335 159 -309
rect 225 -331 255 -309
rect 15 -381 31 -347
rect 65 -381 81 -347
rect 15 -397 81 -381
rect 207 -347 273 -331
rect 321 -335 351 -309
rect 417 -331 447 -309
rect 207 -381 223 -347
rect 257 -381 273 -347
rect 207 -397 273 -381
rect 399 -347 465 -331
rect 399 -381 415 -347
rect 449 -381 465 -347
rect 399 -397 465 -381
rect -369 -455 -303 -439
rect -369 -489 -353 -455
rect -319 -489 -303 -455
rect -447 -527 -417 -501
rect -369 -505 -303 -489
rect -177 -455 -111 -439
rect -177 -489 -161 -455
rect -127 -489 -111 -455
rect -351 -527 -321 -505
rect -255 -527 -225 -501
rect -177 -505 -111 -489
rect 15 -455 81 -439
rect 15 -489 31 -455
rect 65 -489 81 -455
rect -159 -527 -129 -505
rect -63 -527 -33 -501
rect 15 -505 81 -489
rect 207 -455 273 -439
rect 207 -489 223 -455
rect 257 -489 273 -455
rect 33 -527 63 -505
rect 129 -527 159 -501
rect 207 -505 273 -489
rect 399 -455 465 -439
rect 399 -489 415 -455
rect 449 -489 465 -455
rect 225 -527 255 -505
rect 321 -527 351 -501
rect 399 -505 465 -489
rect 417 -527 447 -505
rect -447 -749 -417 -727
rect -465 -765 -399 -749
rect -351 -753 -321 -727
rect -255 -749 -225 -727
rect -465 -799 -449 -765
rect -415 -799 -399 -765
rect -465 -815 -399 -799
rect -273 -765 -207 -749
rect -159 -753 -129 -727
rect -63 -749 -33 -727
rect -273 -799 -257 -765
rect -223 -799 -207 -765
rect -273 -815 -207 -799
rect -81 -765 -15 -749
rect 33 -753 63 -727
rect 129 -749 159 -727
rect -81 -799 -65 -765
rect -31 -799 -15 -765
rect -81 -815 -15 -799
rect 111 -765 177 -749
rect 225 -753 255 -727
rect 321 -749 351 -727
rect 111 -799 127 -765
rect 161 -799 177 -765
rect 111 -815 177 -799
rect 303 -765 369 -749
rect 417 -753 447 -727
rect 303 -799 319 -765
rect 353 -799 369 -765
rect 303 -815 369 -799
<< polycont >>
rect -449 765 -415 799
rect -257 765 -223 799
rect -65 765 -31 799
rect 127 765 161 799
rect 319 765 353 799
rect -353 455 -319 489
rect -161 455 -127 489
rect 31 455 65 489
rect 223 455 257 489
rect 415 455 449 489
rect -353 347 -319 381
rect -161 347 -127 381
rect 31 347 65 381
rect 223 347 257 381
rect 415 347 449 381
rect -449 37 -415 71
rect -257 37 -223 71
rect -65 37 -31 71
rect 127 37 161 71
rect 319 37 353 71
rect -449 -71 -415 -37
rect -257 -71 -223 -37
rect -65 -71 -31 -37
rect 127 -71 161 -37
rect 319 -71 353 -37
rect -353 -381 -319 -347
rect -161 -381 -127 -347
rect 31 -381 65 -347
rect 223 -381 257 -347
rect 415 -381 449 -347
rect -353 -489 -319 -455
rect -161 -489 -127 -455
rect 31 -489 65 -455
rect 223 -489 257 -455
rect 415 -489 449 -455
rect -449 -799 -415 -765
rect -257 -799 -223 -765
rect -65 -799 -31 -765
rect 127 -799 161 -765
rect 319 -799 353 -765
<< locali >>
rect -611 867 -515 901
rect 515 867 611 901
rect -611 805 -577 867
rect 577 805 611 867
rect -465 765 -449 799
rect -415 765 -399 799
rect -273 765 -257 799
rect -223 765 -207 799
rect -81 765 -65 799
rect -31 765 -15 799
rect 111 765 127 799
rect 161 765 177 799
rect 303 765 319 799
rect 353 765 369 799
rect -497 715 -463 731
rect -497 523 -463 539
rect -401 715 -367 731
rect -401 523 -367 539
rect -305 715 -271 731
rect -305 523 -271 539
rect -209 715 -175 731
rect -209 523 -175 539
rect -113 715 -79 731
rect -113 523 -79 539
rect -17 715 17 731
rect -17 523 17 539
rect 79 715 113 731
rect 79 523 113 539
rect 175 715 209 731
rect 175 523 209 539
rect 271 715 305 731
rect 271 523 305 539
rect 367 715 401 731
rect 367 523 401 539
rect 463 715 497 731
rect 463 523 497 539
rect -369 455 -353 489
rect -319 455 -303 489
rect -177 455 -161 489
rect -127 455 -111 489
rect 15 455 31 489
rect 65 455 81 489
rect 207 455 223 489
rect 257 455 273 489
rect 399 455 415 489
rect 449 455 465 489
rect -369 347 -353 381
rect -319 347 -303 381
rect -177 347 -161 381
rect -127 347 -111 381
rect 15 347 31 381
rect 65 347 81 381
rect 207 347 223 381
rect 257 347 273 381
rect 399 347 415 381
rect 449 347 465 381
rect -497 297 -463 313
rect -497 105 -463 121
rect -401 297 -367 313
rect -401 105 -367 121
rect -305 297 -271 313
rect -305 105 -271 121
rect -209 297 -175 313
rect -209 105 -175 121
rect -113 297 -79 313
rect -113 105 -79 121
rect -17 297 17 313
rect -17 105 17 121
rect 79 297 113 313
rect 79 105 113 121
rect 175 297 209 313
rect 175 105 209 121
rect 271 297 305 313
rect 271 105 305 121
rect 367 297 401 313
rect 367 105 401 121
rect 463 297 497 313
rect 463 105 497 121
rect -465 37 -449 71
rect -415 37 -399 71
rect -273 37 -257 71
rect -223 37 -207 71
rect -81 37 -65 71
rect -31 37 -15 71
rect 111 37 127 71
rect 161 37 177 71
rect 303 37 319 71
rect 353 37 369 71
rect -465 -71 -449 -37
rect -415 -71 -399 -37
rect -273 -71 -257 -37
rect -223 -71 -207 -37
rect -81 -71 -65 -37
rect -31 -71 -15 -37
rect 111 -71 127 -37
rect 161 -71 177 -37
rect 303 -71 319 -37
rect 353 -71 369 -37
rect -497 -121 -463 -105
rect -497 -313 -463 -297
rect -401 -121 -367 -105
rect -401 -313 -367 -297
rect -305 -121 -271 -105
rect -305 -313 -271 -297
rect -209 -121 -175 -105
rect -209 -313 -175 -297
rect -113 -121 -79 -105
rect -113 -313 -79 -297
rect -17 -121 17 -105
rect -17 -313 17 -297
rect 79 -121 113 -105
rect 79 -313 113 -297
rect 175 -121 209 -105
rect 175 -313 209 -297
rect 271 -121 305 -105
rect 271 -313 305 -297
rect 367 -121 401 -105
rect 367 -313 401 -297
rect 463 -121 497 -105
rect 463 -313 497 -297
rect -369 -381 -353 -347
rect -319 -381 -303 -347
rect -177 -381 -161 -347
rect -127 -381 -111 -347
rect 15 -381 31 -347
rect 65 -381 81 -347
rect 207 -381 223 -347
rect 257 -381 273 -347
rect 399 -381 415 -347
rect 449 -381 465 -347
rect -369 -489 -353 -455
rect -319 -489 -303 -455
rect -177 -489 -161 -455
rect -127 -489 -111 -455
rect 15 -489 31 -455
rect 65 -489 81 -455
rect 207 -489 223 -455
rect 257 -489 273 -455
rect 399 -489 415 -455
rect 449 -489 465 -455
rect -497 -539 -463 -523
rect -497 -731 -463 -715
rect -401 -539 -367 -523
rect -401 -731 -367 -715
rect -305 -539 -271 -523
rect -305 -731 -271 -715
rect -209 -539 -175 -523
rect -209 -731 -175 -715
rect -113 -539 -79 -523
rect -113 -731 -79 -715
rect -17 -539 17 -523
rect -17 -731 17 -715
rect 79 -539 113 -523
rect 79 -731 113 -715
rect 175 -539 209 -523
rect 175 -731 209 -715
rect 271 -539 305 -523
rect 271 -731 305 -715
rect 367 -539 401 -523
rect 367 -731 401 -715
rect 463 -539 497 -523
rect 463 -731 497 -715
rect -465 -799 -449 -765
rect -415 -799 -399 -765
rect -273 -799 -257 -765
rect -223 -799 -207 -765
rect -81 -799 -65 -765
rect -31 -799 -15 -765
rect 111 -799 127 -765
rect 161 -799 177 -765
rect 303 -799 319 -765
rect 353 -799 369 -765
rect -611 -867 -577 -805
rect 577 -867 611 -805
rect -611 -901 -515 -867
rect 515 -901 611 -867
<< viali >>
rect -449 765 -415 799
rect -257 765 -223 799
rect -65 765 -31 799
rect 127 765 161 799
rect 319 765 353 799
rect -497 539 -463 715
rect -401 539 -367 715
rect -305 539 -271 715
rect -209 539 -175 715
rect -113 539 -79 715
rect -17 539 17 715
rect 79 539 113 715
rect 175 539 209 715
rect 271 539 305 715
rect 367 539 401 715
rect 463 539 497 715
rect -353 455 -319 489
rect -161 455 -127 489
rect 31 455 65 489
rect 223 455 257 489
rect 415 455 449 489
rect -353 347 -319 381
rect -161 347 -127 381
rect 31 347 65 381
rect 223 347 257 381
rect 415 347 449 381
rect -497 121 -463 297
rect -401 121 -367 297
rect -305 121 -271 297
rect -209 121 -175 297
rect -113 121 -79 297
rect -17 121 17 297
rect 79 121 113 297
rect 175 121 209 297
rect 271 121 305 297
rect 367 121 401 297
rect 463 121 497 297
rect -449 37 -415 71
rect -257 37 -223 71
rect -65 37 -31 71
rect 127 37 161 71
rect 319 37 353 71
rect -449 -71 -415 -37
rect -257 -71 -223 -37
rect -65 -71 -31 -37
rect 127 -71 161 -37
rect 319 -71 353 -37
rect -497 -297 -463 -121
rect -401 -297 -367 -121
rect -305 -297 -271 -121
rect -209 -297 -175 -121
rect -113 -297 -79 -121
rect -17 -297 17 -121
rect 79 -297 113 -121
rect 175 -297 209 -121
rect 271 -297 305 -121
rect 367 -297 401 -121
rect 463 -297 497 -121
rect -353 -381 -319 -347
rect -161 -381 -127 -347
rect 31 -381 65 -347
rect 223 -381 257 -347
rect 415 -381 449 -347
rect -353 -489 -319 -455
rect -161 -489 -127 -455
rect 31 -489 65 -455
rect 223 -489 257 -455
rect 415 -489 449 -455
rect -497 -715 -463 -539
rect -401 -715 -367 -539
rect -305 -715 -271 -539
rect -209 -715 -175 -539
rect -113 -715 -79 -539
rect -17 -715 17 -539
rect 79 -715 113 -539
rect 175 -715 209 -539
rect 271 -715 305 -539
rect 367 -715 401 -539
rect 463 -715 497 -539
rect -449 -799 -415 -765
rect -257 -799 -223 -765
rect -65 -799 -31 -765
rect 127 -799 161 -765
rect 319 -799 353 -765
<< metal1 >>
rect -461 799 -403 805
rect -461 765 -449 799
rect -415 765 -403 799
rect -461 759 -403 765
rect -269 799 -211 805
rect -269 765 -257 799
rect -223 765 -211 799
rect -269 759 -211 765
rect -77 799 -19 805
rect -77 765 -65 799
rect -31 765 -19 799
rect -77 759 -19 765
rect 115 799 173 805
rect 115 765 127 799
rect 161 765 173 799
rect 115 759 173 765
rect 307 799 365 805
rect 307 765 319 799
rect 353 765 365 799
rect 307 759 365 765
rect -503 715 -457 727
rect -503 539 -497 715
rect -463 539 -457 715
rect -503 527 -457 539
rect -407 715 -361 727
rect -407 539 -401 715
rect -367 539 -361 715
rect -407 527 -361 539
rect -311 715 -265 727
rect -311 539 -305 715
rect -271 539 -265 715
rect -311 527 -265 539
rect -215 715 -169 727
rect -215 539 -209 715
rect -175 539 -169 715
rect -215 527 -169 539
rect -119 715 -73 727
rect -119 539 -113 715
rect -79 539 -73 715
rect -119 527 -73 539
rect -23 715 23 727
rect -23 539 -17 715
rect 17 539 23 715
rect -23 527 23 539
rect 73 715 119 727
rect 73 539 79 715
rect 113 539 119 715
rect 73 527 119 539
rect 169 715 215 727
rect 169 539 175 715
rect 209 539 215 715
rect 169 527 215 539
rect 265 715 311 727
rect 265 539 271 715
rect 305 539 311 715
rect 265 527 311 539
rect 361 715 407 727
rect 361 539 367 715
rect 401 539 407 715
rect 361 527 407 539
rect 457 715 503 727
rect 457 539 463 715
rect 497 539 503 715
rect 457 527 503 539
rect -365 489 -307 495
rect -365 455 -353 489
rect -319 455 -307 489
rect -365 449 -307 455
rect -173 489 -115 495
rect -173 455 -161 489
rect -127 455 -115 489
rect -173 449 -115 455
rect 19 489 77 495
rect 19 455 31 489
rect 65 455 77 489
rect 19 449 77 455
rect 211 489 269 495
rect 211 455 223 489
rect 257 455 269 489
rect 211 449 269 455
rect 403 489 461 495
rect 403 455 415 489
rect 449 455 461 489
rect 403 449 461 455
rect -365 381 -307 387
rect -365 347 -353 381
rect -319 347 -307 381
rect -365 341 -307 347
rect -173 381 -115 387
rect -173 347 -161 381
rect -127 347 -115 381
rect -173 341 -115 347
rect 19 381 77 387
rect 19 347 31 381
rect 65 347 77 381
rect 19 341 77 347
rect 211 381 269 387
rect 211 347 223 381
rect 257 347 269 381
rect 211 341 269 347
rect 403 381 461 387
rect 403 347 415 381
rect 449 347 461 381
rect 403 341 461 347
rect -503 297 -457 309
rect -503 121 -497 297
rect -463 121 -457 297
rect -503 109 -457 121
rect -407 297 -361 309
rect -407 121 -401 297
rect -367 121 -361 297
rect -407 109 -361 121
rect -311 297 -265 309
rect -311 121 -305 297
rect -271 121 -265 297
rect -311 109 -265 121
rect -215 297 -169 309
rect -215 121 -209 297
rect -175 121 -169 297
rect -215 109 -169 121
rect -119 297 -73 309
rect -119 121 -113 297
rect -79 121 -73 297
rect -119 109 -73 121
rect -23 297 23 309
rect -23 121 -17 297
rect 17 121 23 297
rect -23 109 23 121
rect 73 297 119 309
rect 73 121 79 297
rect 113 121 119 297
rect 73 109 119 121
rect 169 297 215 309
rect 169 121 175 297
rect 209 121 215 297
rect 169 109 215 121
rect 265 297 311 309
rect 265 121 271 297
rect 305 121 311 297
rect 265 109 311 121
rect 361 297 407 309
rect 361 121 367 297
rect 401 121 407 297
rect 361 109 407 121
rect 457 297 503 309
rect 457 121 463 297
rect 497 121 503 297
rect 457 109 503 121
rect -461 71 -403 77
rect -461 37 -449 71
rect -415 37 -403 71
rect -461 31 -403 37
rect -269 71 -211 77
rect -269 37 -257 71
rect -223 37 -211 71
rect -269 31 -211 37
rect -77 71 -19 77
rect -77 37 -65 71
rect -31 37 -19 71
rect -77 31 -19 37
rect 115 71 173 77
rect 115 37 127 71
rect 161 37 173 71
rect 115 31 173 37
rect 307 71 365 77
rect 307 37 319 71
rect 353 37 365 71
rect 307 31 365 37
rect -461 -37 -403 -31
rect -461 -71 -449 -37
rect -415 -71 -403 -37
rect -461 -77 -403 -71
rect -269 -37 -211 -31
rect -269 -71 -257 -37
rect -223 -71 -211 -37
rect -269 -77 -211 -71
rect -77 -37 -19 -31
rect -77 -71 -65 -37
rect -31 -71 -19 -37
rect -77 -77 -19 -71
rect 115 -37 173 -31
rect 115 -71 127 -37
rect 161 -71 173 -37
rect 115 -77 173 -71
rect 307 -37 365 -31
rect 307 -71 319 -37
rect 353 -71 365 -37
rect 307 -77 365 -71
rect -503 -121 -457 -109
rect -503 -297 -497 -121
rect -463 -297 -457 -121
rect -503 -309 -457 -297
rect -407 -121 -361 -109
rect -407 -297 -401 -121
rect -367 -297 -361 -121
rect -407 -309 -361 -297
rect -311 -121 -265 -109
rect -311 -297 -305 -121
rect -271 -297 -265 -121
rect -311 -309 -265 -297
rect -215 -121 -169 -109
rect -215 -297 -209 -121
rect -175 -297 -169 -121
rect -215 -309 -169 -297
rect -119 -121 -73 -109
rect -119 -297 -113 -121
rect -79 -297 -73 -121
rect -119 -309 -73 -297
rect -23 -121 23 -109
rect -23 -297 -17 -121
rect 17 -297 23 -121
rect -23 -309 23 -297
rect 73 -121 119 -109
rect 73 -297 79 -121
rect 113 -297 119 -121
rect 73 -309 119 -297
rect 169 -121 215 -109
rect 169 -297 175 -121
rect 209 -297 215 -121
rect 169 -309 215 -297
rect 265 -121 311 -109
rect 265 -297 271 -121
rect 305 -297 311 -121
rect 265 -309 311 -297
rect 361 -121 407 -109
rect 361 -297 367 -121
rect 401 -297 407 -121
rect 361 -309 407 -297
rect 457 -121 503 -109
rect 457 -297 463 -121
rect 497 -297 503 -121
rect 457 -309 503 -297
rect -365 -347 -307 -341
rect -365 -381 -353 -347
rect -319 -381 -307 -347
rect -365 -387 -307 -381
rect -173 -347 -115 -341
rect -173 -381 -161 -347
rect -127 -381 -115 -347
rect -173 -387 -115 -381
rect 19 -347 77 -341
rect 19 -381 31 -347
rect 65 -381 77 -347
rect 19 -387 77 -381
rect 211 -347 269 -341
rect 211 -381 223 -347
rect 257 -381 269 -347
rect 211 -387 269 -381
rect 403 -347 461 -341
rect 403 -381 415 -347
rect 449 -381 461 -347
rect 403 -387 461 -381
rect -365 -455 -307 -449
rect -365 -489 -353 -455
rect -319 -489 -307 -455
rect -365 -495 -307 -489
rect -173 -455 -115 -449
rect -173 -489 -161 -455
rect -127 -489 -115 -455
rect -173 -495 -115 -489
rect 19 -455 77 -449
rect 19 -489 31 -455
rect 65 -489 77 -455
rect 19 -495 77 -489
rect 211 -455 269 -449
rect 211 -489 223 -455
rect 257 -489 269 -455
rect 211 -495 269 -489
rect 403 -455 461 -449
rect 403 -489 415 -455
rect 449 -489 461 -455
rect 403 -495 461 -489
rect -503 -539 -457 -527
rect -503 -715 -497 -539
rect -463 -715 -457 -539
rect -503 -727 -457 -715
rect -407 -539 -361 -527
rect -407 -715 -401 -539
rect -367 -715 -361 -539
rect -407 -727 -361 -715
rect -311 -539 -265 -527
rect -311 -715 -305 -539
rect -271 -715 -265 -539
rect -311 -727 -265 -715
rect -215 -539 -169 -527
rect -215 -715 -209 -539
rect -175 -715 -169 -539
rect -215 -727 -169 -715
rect -119 -539 -73 -527
rect -119 -715 -113 -539
rect -79 -715 -73 -539
rect -119 -727 -73 -715
rect -23 -539 23 -527
rect -23 -715 -17 -539
rect 17 -715 23 -539
rect -23 -727 23 -715
rect 73 -539 119 -527
rect 73 -715 79 -539
rect 113 -715 119 -539
rect 73 -727 119 -715
rect 169 -539 215 -527
rect 169 -715 175 -539
rect 209 -715 215 -539
rect 169 -727 215 -715
rect 265 -539 311 -527
rect 265 -715 271 -539
rect 305 -715 311 -539
rect 265 -727 311 -715
rect 361 -539 407 -527
rect 361 -715 367 -539
rect 401 -715 407 -539
rect 361 -727 407 -715
rect 457 -539 503 -527
rect 457 -715 463 -539
rect 497 -715 503 -539
rect 457 -727 503 -715
rect -461 -765 -403 -759
rect -461 -799 -449 -765
rect -415 -799 -403 -765
rect -461 -805 -403 -799
rect -269 -765 -211 -759
rect -269 -799 -257 -765
rect -223 -799 -211 -765
rect -269 -805 -211 -799
rect -77 -765 -19 -759
rect -77 -799 -65 -765
rect -31 -799 -19 -765
rect -77 -805 -19 -799
rect 115 -765 173 -759
rect 115 -799 127 -765
rect 161 -799 173 -765
rect 115 -805 173 -799
rect 307 -765 365 -759
rect 307 -799 319 -765
rect 353 -799 365 -765
rect 307 -805 365 -799
<< properties >>
string FIXED_BBOX -594 -884 594 884
string gencell sky130_fd_pr__nfet_01v8_lvt
string library sky130
string parameters w 1.0 l 0.15 m 4 nf 10 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
