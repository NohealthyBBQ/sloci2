magic
tech sky130A
magscale 1 2
timestamp 1672462443
<< dnwell >>
rect -1960 1360 1960 1960
rect -1960 -1360 -1360 1360
rect 1360 -1360 1960 1360
rect -1960 -1960 1960 -1360
<< photodiode >>
rect -300 -300 300 300
<< nwell >>
rect -2040 1754 2040 2040
rect -2040 -1754 -1754 1754
rect -84 -84 84 84
rect 1754 -1754 2040 1754
rect -2040 -2040 2040 -1754
<< pwell >>
rect -2147 2041 2147 2147
rect -2147 -2041 -2041 2041
rect 2041 -2041 2147 2041
rect -2147 -2147 2147 -2041
<< psubdiff >>
rect -2111 2077 -2015 2111
rect 2015 2077 2111 2111
rect -2111 2015 -2077 2077
rect 2077 2015 2111 2077
rect -2111 -2077 -2077 -2015
rect 2077 -2077 2111 -2015
rect -2111 -2111 -2015 -2077
rect 2015 -2111 2111 -2077
<< nsubdiff >>
rect -1914 1880 -1818 1914
rect 1818 1880 1914 1914
rect -1914 1818 -1880 1880
rect 1880 1818 1914 1880
rect -41 17 41 41
rect -41 -17 -17 17
rect 17 -17 41 17
rect -41 -41 41 -17
rect -1914 -1880 -1880 -1818
rect 1880 -1880 1914 -1818
rect -1914 -1914 -1818 -1880
rect 1818 -1914 1914 -1880
<< psubdiffcont >>
rect -2015 2077 2015 2111
rect -2111 -2015 -2077 2015
rect 2077 -2015 2111 2015
rect -2015 -2111 2015 -2077
<< nsubdiffcont >>
rect -1818 1880 1818 1914
rect -1914 -1818 -1880 1818
rect -17 -17 17 17
rect 1880 -1818 1914 1818
rect -1818 -1914 1818 -1880
<< locali >>
rect -2111 2077 -2015 2111
rect 2015 2077 2111 2111
rect -2111 2015 -2077 2077
rect 2077 2015 2111 2077
rect -1914 1880 -1818 1914
rect 1818 1880 1914 1914
rect -1914 1818 -1880 1880
rect 1880 1818 1914 1880
rect -33 -17 -17 17
rect 17 -17 33 17
rect -1914 -1880 -1880 -1818
rect 1880 -1880 1914 -1818
rect -1914 -1914 -1818 -1880
rect 1818 -1914 1914 -1880
rect -2111 -2077 -2077 -2015
rect 2077 -2077 2111 -2015
rect -2111 -2111 -2015 -2077
rect 2015 -2111 2111 -2077
<< properties >>
string FIXED_BBOX -2094 -2094 2094 2094
string gencell sky130_fd_pr__photodiode
string library sky130
string parameters nx 1 ny 1 deltax 0 deltay 0 xstep 8.0 ystep 8.0
<< end >>
