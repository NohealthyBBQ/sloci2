magic
tech sky130A
magscale 1 2
timestamp 1662826682
<< pwell >>
rect -739 -55534 739 55534
<< psubdiff >>
rect -703 55464 -607 55498
rect 607 55464 703 55498
rect -703 55402 -669 55464
rect 669 55402 703 55464
rect -703 -55464 -669 -55402
rect 669 -55464 703 -55402
rect -703 -55498 -607 -55464
rect 607 -55498 703 -55464
<< psubdiffcont >>
rect -607 55464 607 55498
rect -703 -55402 -669 55402
rect 669 -55402 703 55402
rect -607 -55498 607 -55464
<< xpolycontact >>
rect -573 54936 573 55368
rect -573 33304 573 33736
rect -573 32768 573 33200
rect -573 11136 573 11568
rect -573 10600 573 11032
rect -573 -11032 573 -10600
rect -573 -11568 573 -11136
rect -573 -33200 573 -32768
rect -573 -33736 573 -33304
rect -573 -55368 573 -54936
<< xpolyres >>
rect -573 33736 573 54936
rect -573 11568 573 32768
rect -573 -10600 573 10600
rect -573 -32768 573 -11568
rect -573 -54936 573 -33736
<< locali >>
rect -703 55464 -607 55498
rect 607 55464 703 55498
rect -703 55402 -669 55464
rect 669 55402 703 55464
rect -703 -55464 -669 -55402
rect 669 -55464 703 -55402
rect -703 -55498 -607 -55464
rect 607 -55498 703 -55464
<< viali >>
rect -557 54953 557 55350
rect -557 33322 557 33719
rect -557 32785 557 33182
rect -557 11154 557 11551
rect -557 10617 557 11014
rect -557 -11014 557 -10617
rect -557 -11551 557 -11154
rect -557 -33182 557 -32785
rect -557 -33719 557 -33322
rect -557 -55350 557 -54953
<< metal1 >>
rect -569 55350 569 55356
rect -569 54953 -557 55350
rect 557 54953 569 55350
rect -569 54947 569 54953
rect -569 33719 569 33725
rect -569 33322 -557 33719
rect 557 33322 569 33719
rect -569 33316 569 33322
rect -569 33182 569 33188
rect -569 32785 -557 33182
rect 557 32785 569 33182
rect -569 32779 569 32785
rect -569 11551 569 11557
rect -569 11154 -557 11551
rect 557 11154 569 11551
rect -569 11148 569 11154
rect -569 11014 569 11020
rect -569 10617 -557 11014
rect 557 10617 569 11014
rect -569 10611 569 10617
rect -569 -10617 569 -10611
rect -569 -11014 -557 -10617
rect 557 -11014 569 -10617
rect -569 -11020 569 -11014
rect -569 -11154 569 -11148
rect -569 -11551 -557 -11154
rect 557 -11551 569 -11154
rect -569 -11557 569 -11551
rect -569 -32785 569 -32779
rect -569 -33182 -557 -32785
rect 557 -33182 569 -32785
rect -569 -33188 569 -33182
rect -569 -33322 569 -33316
rect -569 -33719 -557 -33322
rect 557 -33719 569 -33322
rect -569 -33725 569 -33719
rect -569 -54953 569 -54947
rect -569 -55350 -557 -54953
rect 557 -55350 569 -54953
rect -569 -55356 569 -55350
<< res5p73 >>
rect -575 33734 575 54938
rect -575 11566 575 32770
rect -575 -10602 575 10602
rect -575 -32770 575 -11566
rect -575 -54938 575 -33734
<< properties >>
string FIXED_BBOX -686 -55481 686 55481
string gencell sky130_fd_pr__res_xhigh_po_5p73
string library sky130
string parameters w 5.730 l 106 m 5 nx 1 wmin 5.730 lmin 0.50 rho 2000 val 37.063k dummy 0 dw 0.0 term 188.2 sterm 0.0 caplen 0 wmax 5.730 guard 1 glc 1 grc 1 gtc 1 gbc 1 compatible {sky130_fd_pr__res_xhigh_po_0p35  sky130_fd_pr__res_xhigh_po_0p69 sky130_fd_pr__res_xhigh_po_1p41  sky130_fd_pr__res_xhigh_po_2p85 sky130_fd_pr__res_xhigh_po_5p73} snake 0 full_metal 1 n_guard 0 hv_guard 0 vias 1 viagb 0 viagt 0 viagl 0 viagr 0
<< end >>
