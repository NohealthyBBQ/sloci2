magic
tech sky130A
magscale 1 2
timestamp 1672484988
<< metal1 >>
rect 5046 2024 5108 2106
rect 5122 1930 5390 1974
rect 5380 1922 5390 1930
rect 5442 1922 5452 1974
rect 4950 1856 5040 1884
rect 4950 1758 4978 1856
rect 4912 1702 4922 1758
rect 4978 1702 4988 1758
rect 5022 1714 5134 1748
rect 4950 1598 4960 1650
rect 5012 1598 5022 1650
rect 5136 1478 5160 1530
rect 5212 1478 5222 1530
rect 5136 1472 5212 1478
rect 5046 1352 5108 1434
<< via1 >>
rect 5390 1922 5442 1974
rect 4922 1702 4978 1758
rect 4960 1598 5012 1650
rect 5160 1478 5212 1530
<< metal2 >>
rect 5390 1974 5442 1984
rect 4806 1624 4834 1952
rect 5390 1912 5442 1922
rect 4922 1758 4978 1768
rect 4922 1692 4978 1702
rect 4960 1650 5012 1660
rect 4806 1598 4960 1624
rect 4806 1592 5012 1598
rect 4960 1588 5012 1592
rect 5160 1530 5212 1540
rect 5160 1468 5212 1478
<< via2 >>
rect 4922 1702 4978 1758
<< metal3 >>
rect 4930 1763 5604 1764
rect 4912 1758 5604 1763
rect 4912 1702 4922 1758
rect 4978 1702 5604 1758
rect 4912 1697 4988 1702
use cons1  cons1_0
timestamp 1672483164
transform 1 0 -46340 0 1 8198
box 46340 -8198 69992 -4736
use sky130_fd_pr__nfet_01v8_lvt_595QY5  sky130_fd_pr__nfet_01v8_lvt_595QY5_0
timestamp 1672483605
transform 1 0 5077 0 1 1576
box -73 -188 73 188
use sky130_fd_pr__nfet_01v8_lvt_595QY5  sky130_fd_pr__nfet_01v8_lvt_595QY5_1
timestamp 1672483605
transform 1 0 5077 0 1 1886
box -73 -188 73 188
<< end >>
