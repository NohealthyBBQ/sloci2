magic
tech sky130A
magscale 1 2
timestamp 1661905147
<< pwell >>
rect -1312 -657 1312 657
<< nmoslvt >>
rect -1116 109 -716 509
rect -658 109 -258 509
rect -200 109 200 509
rect 258 109 658 509
rect 716 109 1116 509
rect -1116 -447 -716 -47
rect -658 -447 -258 -47
rect -200 -447 200 -47
rect 258 -447 658 -47
rect 716 -447 1116 -47
<< ndiff >>
rect -1174 497 -1116 509
rect -1174 121 -1162 497
rect -1128 121 -1116 497
rect -1174 109 -1116 121
rect -716 497 -658 509
rect -716 121 -704 497
rect -670 121 -658 497
rect -716 109 -658 121
rect -258 497 -200 509
rect -258 121 -246 497
rect -212 121 -200 497
rect -258 109 -200 121
rect 200 497 258 509
rect 200 121 212 497
rect 246 121 258 497
rect 200 109 258 121
rect 658 497 716 509
rect 658 121 670 497
rect 704 121 716 497
rect 658 109 716 121
rect 1116 497 1174 509
rect 1116 121 1128 497
rect 1162 121 1174 497
rect 1116 109 1174 121
rect -1174 -59 -1116 -47
rect -1174 -435 -1162 -59
rect -1128 -435 -1116 -59
rect -1174 -447 -1116 -435
rect -716 -59 -658 -47
rect -716 -435 -704 -59
rect -670 -435 -658 -59
rect -716 -447 -658 -435
rect -258 -59 -200 -47
rect -258 -435 -246 -59
rect -212 -435 -200 -59
rect -258 -447 -200 -435
rect 200 -59 258 -47
rect 200 -435 212 -59
rect 246 -435 258 -59
rect 200 -447 258 -435
rect 658 -59 716 -47
rect 658 -435 670 -59
rect 704 -435 716 -59
rect 658 -447 716 -435
rect 1116 -59 1174 -47
rect 1116 -435 1128 -59
rect 1162 -435 1174 -59
rect 1116 -447 1174 -435
<< ndiffc >>
rect -1162 121 -1128 497
rect -704 121 -670 497
rect -246 121 -212 497
rect 212 121 246 497
rect 670 121 704 497
rect 1128 121 1162 497
rect -1162 -435 -1128 -59
rect -704 -435 -670 -59
rect -246 -435 -212 -59
rect 212 -435 246 -59
rect 670 -435 704 -59
rect 1128 -435 1162 -59
<< psubdiff >>
rect -1276 587 -1180 621
rect 1180 587 1276 621
rect -1276 525 -1242 587
rect 1242 525 1276 587
rect -1276 -587 -1242 -525
rect 1242 -587 1276 -525
rect -1276 -621 -1180 -587
rect 1180 -621 1276 -587
<< psubdiffcont >>
rect -1180 587 1180 621
rect -1276 -525 -1242 525
rect 1242 -525 1276 525
rect -1180 -621 1180 -587
<< poly >>
rect -1116 509 -716 535
rect -658 509 -258 535
rect -200 509 200 535
rect 258 509 658 535
rect 716 509 1116 535
rect -1116 71 -716 109
rect -1116 37 -1100 71
rect -732 37 -716 71
rect -1116 21 -716 37
rect -658 71 -258 109
rect -658 37 -642 71
rect -274 37 -258 71
rect -658 21 -258 37
rect -200 71 200 109
rect -200 37 -184 71
rect 184 37 200 71
rect -200 21 200 37
rect 258 71 658 109
rect 258 37 274 71
rect 642 37 658 71
rect 258 21 658 37
rect 716 71 1116 109
rect 716 37 732 71
rect 1100 37 1116 71
rect 716 21 1116 37
rect -1116 -47 -716 -21
rect -658 -47 -258 -21
rect -200 -47 200 -21
rect 258 -47 658 -21
rect 716 -47 1116 -21
rect -1116 -485 -716 -447
rect -1116 -519 -1100 -485
rect -732 -519 -716 -485
rect -1116 -535 -716 -519
rect -658 -485 -258 -447
rect -658 -519 -642 -485
rect -274 -519 -258 -485
rect -658 -535 -258 -519
rect -200 -485 200 -447
rect -200 -519 -184 -485
rect 184 -519 200 -485
rect -200 -535 200 -519
rect 258 -485 658 -447
rect 258 -519 274 -485
rect 642 -519 658 -485
rect 258 -535 658 -519
rect 716 -485 1116 -447
rect 716 -519 732 -485
rect 1100 -519 1116 -485
rect 716 -535 1116 -519
<< polycont >>
rect -1100 37 -732 71
rect -642 37 -274 71
rect -184 37 184 71
rect 274 37 642 71
rect 732 37 1100 71
rect -1100 -519 -732 -485
rect -642 -519 -274 -485
rect -184 -519 184 -485
rect 274 -519 642 -485
rect 732 -519 1100 -485
<< locali >>
rect -1276 587 -1180 621
rect 1180 587 1276 621
rect -1276 525 -1242 587
rect 1242 525 1276 587
rect -1162 497 -1128 513
rect -1162 105 -1128 121
rect -704 497 -670 513
rect -704 105 -670 121
rect -246 497 -212 513
rect -246 105 -212 121
rect 212 497 246 513
rect 212 105 246 121
rect 670 497 704 513
rect 670 105 704 121
rect 1128 497 1162 513
rect 1128 105 1162 121
rect -1116 37 -1100 71
rect -732 37 -716 71
rect -658 37 -642 71
rect -274 37 -258 71
rect -200 37 -184 71
rect 184 37 200 71
rect 258 37 274 71
rect 642 37 658 71
rect 716 37 732 71
rect 1100 37 1116 71
rect -1162 -59 -1128 -43
rect -1162 -451 -1128 -435
rect -704 -59 -670 -43
rect -704 -451 -670 -435
rect -246 -59 -212 -43
rect -246 -451 -212 -435
rect 212 -59 246 -43
rect 212 -451 246 -435
rect 670 -59 704 -43
rect 670 -451 704 -435
rect 1128 -59 1162 -43
rect 1128 -451 1162 -435
rect -1116 -519 -1100 -485
rect -732 -519 -716 -485
rect -658 -519 -642 -485
rect -274 -519 -258 -485
rect -200 -519 -184 -485
rect 184 -519 200 -485
rect 258 -519 274 -485
rect 642 -519 658 -485
rect 716 -519 732 -485
rect 1100 -519 1116 -485
rect -1276 -587 -1242 -525
rect 1242 -587 1276 -525
rect -1276 -621 -1180 -587
rect 1180 -621 1276 -587
<< viali >>
rect -1162 121 -1128 497
rect -704 121 -670 497
rect -246 121 -212 497
rect 212 121 246 497
rect 670 121 704 497
rect 1128 121 1162 497
rect -1100 37 -732 71
rect -642 37 -274 71
rect -184 37 184 71
rect 274 37 642 71
rect 732 37 1100 71
rect -1162 -435 -1128 -59
rect -704 -435 -670 -59
rect -246 -435 -212 -59
rect 212 -435 246 -59
rect 670 -435 704 -59
rect 1128 -435 1162 -59
rect -1100 -519 -732 -485
rect -642 -519 -274 -485
rect -184 -519 184 -485
rect 274 -519 642 -485
rect 732 -519 1100 -485
<< metal1 >>
rect -1168 497 -1122 509
rect -1168 121 -1162 497
rect -1128 121 -1122 497
rect -1168 109 -1122 121
rect -710 497 -664 509
rect -710 121 -704 497
rect -670 121 -664 497
rect -710 109 -664 121
rect -252 497 -206 509
rect -252 121 -246 497
rect -212 121 -206 497
rect -252 109 -206 121
rect 206 497 252 509
rect 206 121 212 497
rect 246 121 252 497
rect 206 109 252 121
rect 664 497 710 509
rect 664 121 670 497
rect 704 121 710 497
rect 664 109 710 121
rect 1122 497 1168 509
rect 1122 121 1128 497
rect 1162 121 1168 497
rect 1122 109 1168 121
rect -1112 71 -720 77
rect -1112 37 -1100 71
rect -732 37 -720 71
rect -1112 31 -720 37
rect -654 71 -262 77
rect -654 37 -642 71
rect -274 37 -262 71
rect -654 31 -262 37
rect -196 71 196 77
rect -196 37 -184 71
rect 184 37 196 71
rect -196 31 196 37
rect 262 71 654 77
rect 262 37 274 71
rect 642 37 654 71
rect 262 31 654 37
rect 720 71 1112 77
rect 720 37 732 71
rect 1100 37 1112 71
rect 720 31 1112 37
rect -1168 -59 -1122 -47
rect -1168 -435 -1162 -59
rect -1128 -435 -1122 -59
rect -1168 -447 -1122 -435
rect -710 -59 -664 -47
rect -710 -435 -704 -59
rect -670 -435 -664 -59
rect -710 -447 -664 -435
rect -252 -59 -206 -47
rect -252 -435 -246 -59
rect -212 -435 -206 -59
rect -252 -447 -206 -435
rect 206 -59 252 -47
rect 206 -435 212 -59
rect 246 -435 252 -59
rect 206 -447 252 -435
rect 664 -59 710 -47
rect 664 -435 670 -59
rect 704 -435 710 -59
rect 664 -447 710 -435
rect 1122 -59 1168 -47
rect 1122 -435 1128 -59
rect 1162 -435 1168 -59
rect 1122 -447 1168 -435
rect -1112 -485 -720 -479
rect -1112 -519 -1100 -485
rect -732 -519 -720 -485
rect -1112 -525 -720 -519
rect -654 -485 -262 -479
rect -654 -519 -642 -485
rect -274 -519 -262 -485
rect -654 -525 -262 -519
rect -196 -485 196 -479
rect -196 -519 -184 -485
rect 184 -519 196 -485
rect -196 -525 196 -519
rect 262 -485 654 -479
rect 262 -519 274 -485
rect 642 -519 654 -485
rect 262 -525 654 -519
rect 720 -485 1112 -479
rect 720 -519 732 -485
rect 1100 -519 1112 -485
rect 720 -525 1112 -519
<< properties >>
string FIXED_BBOX -1259 -604 1259 604
string gencell sky130_fd_pr__nfet_01v8_lvt
string library sky130
string parameters w 2 l 2 m 2 nf 5 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 0 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
