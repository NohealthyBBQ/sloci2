magic
tech sky130A
magscale 1 2
timestamp 1672264357
<< nwell >>
rect -2686 -3537 2686 3537
<< pmoslvt >>
rect -2490 118 -2090 3318
rect -2032 118 -1632 3318
rect -1574 118 -1174 3318
rect -1116 118 -716 3318
rect -658 118 -258 3318
rect -200 118 200 3318
rect 258 118 658 3318
rect 716 118 1116 3318
rect 1174 118 1574 3318
rect 1632 118 2032 3318
rect 2090 118 2490 3318
rect -2490 -3318 -2090 -118
rect -2032 -3318 -1632 -118
rect -1574 -3318 -1174 -118
rect -1116 -3318 -716 -118
rect -658 -3318 -258 -118
rect -200 -3318 200 -118
rect 258 -3318 658 -118
rect 716 -3318 1116 -118
rect 1174 -3318 1574 -118
rect 1632 -3318 2032 -118
rect 2090 -3318 2490 -118
<< pdiff >>
rect -2548 3306 -2490 3318
rect -2548 130 -2536 3306
rect -2502 130 -2490 3306
rect -2548 118 -2490 130
rect -2090 3306 -2032 3318
rect -2090 130 -2078 3306
rect -2044 130 -2032 3306
rect -2090 118 -2032 130
rect -1632 3306 -1574 3318
rect -1632 130 -1620 3306
rect -1586 130 -1574 3306
rect -1632 118 -1574 130
rect -1174 3306 -1116 3318
rect -1174 130 -1162 3306
rect -1128 130 -1116 3306
rect -1174 118 -1116 130
rect -716 3306 -658 3318
rect -716 130 -704 3306
rect -670 130 -658 3306
rect -716 118 -658 130
rect -258 3306 -200 3318
rect -258 130 -246 3306
rect -212 130 -200 3306
rect -258 118 -200 130
rect 200 3306 258 3318
rect 200 130 212 3306
rect 246 130 258 3306
rect 200 118 258 130
rect 658 3306 716 3318
rect 658 130 670 3306
rect 704 130 716 3306
rect 658 118 716 130
rect 1116 3306 1174 3318
rect 1116 130 1128 3306
rect 1162 130 1174 3306
rect 1116 118 1174 130
rect 1574 3306 1632 3318
rect 1574 130 1586 3306
rect 1620 130 1632 3306
rect 1574 118 1632 130
rect 2032 3306 2090 3318
rect 2032 130 2044 3306
rect 2078 130 2090 3306
rect 2032 118 2090 130
rect 2490 3306 2548 3318
rect 2490 130 2502 3306
rect 2536 130 2548 3306
rect 2490 118 2548 130
rect -2548 -130 -2490 -118
rect -2548 -3306 -2536 -130
rect -2502 -3306 -2490 -130
rect -2548 -3318 -2490 -3306
rect -2090 -130 -2032 -118
rect -2090 -3306 -2078 -130
rect -2044 -3306 -2032 -130
rect -2090 -3318 -2032 -3306
rect -1632 -130 -1574 -118
rect -1632 -3306 -1620 -130
rect -1586 -3306 -1574 -130
rect -1632 -3318 -1574 -3306
rect -1174 -130 -1116 -118
rect -1174 -3306 -1162 -130
rect -1128 -3306 -1116 -130
rect -1174 -3318 -1116 -3306
rect -716 -130 -658 -118
rect -716 -3306 -704 -130
rect -670 -3306 -658 -130
rect -716 -3318 -658 -3306
rect -258 -130 -200 -118
rect -258 -3306 -246 -130
rect -212 -3306 -200 -130
rect -258 -3318 -200 -3306
rect 200 -130 258 -118
rect 200 -3306 212 -130
rect 246 -3306 258 -130
rect 200 -3318 258 -3306
rect 658 -130 716 -118
rect 658 -3306 670 -130
rect 704 -3306 716 -130
rect 658 -3318 716 -3306
rect 1116 -130 1174 -118
rect 1116 -3306 1128 -130
rect 1162 -3306 1174 -130
rect 1116 -3318 1174 -3306
rect 1574 -130 1632 -118
rect 1574 -3306 1586 -130
rect 1620 -3306 1632 -130
rect 1574 -3318 1632 -3306
rect 2032 -130 2090 -118
rect 2032 -3306 2044 -130
rect 2078 -3306 2090 -130
rect 2032 -3318 2090 -3306
rect 2490 -130 2548 -118
rect 2490 -3306 2502 -130
rect 2536 -3306 2548 -130
rect 2490 -3318 2548 -3306
<< pdiffc >>
rect -2536 130 -2502 3306
rect -2078 130 -2044 3306
rect -1620 130 -1586 3306
rect -1162 130 -1128 3306
rect -704 130 -670 3306
rect -246 130 -212 3306
rect 212 130 246 3306
rect 670 130 704 3306
rect 1128 130 1162 3306
rect 1586 130 1620 3306
rect 2044 130 2078 3306
rect 2502 130 2536 3306
rect -2536 -3306 -2502 -130
rect -2078 -3306 -2044 -130
rect -1620 -3306 -1586 -130
rect -1162 -3306 -1128 -130
rect -704 -3306 -670 -130
rect -246 -3306 -212 -130
rect 212 -3306 246 -130
rect 670 -3306 704 -130
rect 1128 -3306 1162 -130
rect 1586 -3306 1620 -130
rect 2044 -3306 2078 -130
rect 2502 -3306 2536 -130
<< nsubdiff >>
rect -2650 3467 -2554 3501
rect 2554 3467 2650 3501
rect -2650 3405 -2616 3467
rect 2616 3405 2650 3467
rect -2650 -3467 -2616 -3405
rect 2616 -3467 2650 -3405
rect -2650 -3501 -2554 -3467
rect 2554 -3501 2650 -3467
<< nsubdiffcont >>
rect -2554 3467 2554 3501
rect -2650 -3405 -2616 3405
rect 2616 -3405 2650 3405
rect -2554 -3501 2554 -3467
<< poly >>
rect -2490 3399 -2090 3415
rect -2490 3365 -2474 3399
rect -2106 3365 -2090 3399
rect -2490 3318 -2090 3365
rect -2032 3399 -1632 3415
rect -2032 3365 -2016 3399
rect -1648 3365 -1632 3399
rect -2032 3318 -1632 3365
rect -1574 3399 -1174 3415
rect -1574 3365 -1558 3399
rect -1190 3365 -1174 3399
rect -1574 3318 -1174 3365
rect -1116 3399 -716 3415
rect -1116 3365 -1100 3399
rect -732 3365 -716 3399
rect -1116 3318 -716 3365
rect -658 3399 -258 3415
rect -658 3365 -642 3399
rect -274 3365 -258 3399
rect -658 3318 -258 3365
rect -200 3399 200 3415
rect -200 3365 -184 3399
rect 184 3365 200 3399
rect -200 3318 200 3365
rect 258 3399 658 3415
rect 258 3365 274 3399
rect 642 3365 658 3399
rect 258 3318 658 3365
rect 716 3399 1116 3415
rect 716 3365 732 3399
rect 1100 3365 1116 3399
rect 716 3318 1116 3365
rect 1174 3399 1574 3415
rect 1174 3365 1190 3399
rect 1558 3365 1574 3399
rect 1174 3318 1574 3365
rect 1632 3399 2032 3415
rect 1632 3365 1648 3399
rect 2016 3365 2032 3399
rect 1632 3318 2032 3365
rect 2090 3399 2490 3415
rect 2090 3365 2106 3399
rect 2474 3365 2490 3399
rect 2090 3318 2490 3365
rect -2490 71 -2090 118
rect -2490 37 -2474 71
rect -2106 37 -2090 71
rect -2490 21 -2090 37
rect -2032 71 -1632 118
rect -2032 37 -2016 71
rect -1648 37 -1632 71
rect -2032 21 -1632 37
rect -1574 71 -1174 118
rect -1574 37 -1558 71
rect -1190 37 -1174 71
rect -1574 21 -1174 37
rect -1116 71 -716 118
rect -1116 37 -1100 71
rect -732 37 -716 71
rect -1116 21 -716 37
rect -658 71 -258 118
rect -658 37 -642 71
rect -274 37 -258 71
rect -658 21 -258 37
rect -200 71 200 118
rect -200 37 -184 71
rect 184 37 200 71
rect -200 21 200 37
rect 258 71 658 118
rect 258 37 274 71
rect 642 37 658 71
rect 258 21 658 37
rect 716 71 1116 118
rect 716 37 732 71
rect 1100 37 1116 71
rect 716 21 1116 37
rect 1174 71 1574 118
rect 1174 37 1190 71
rect 1558 37 1574 71
rect 1174 21 1574 37
rect 1632 71 2032 118
rect 1632 37 1648 71
rect 2016 37 2032 71
rect 1632 21 2032 37
rect 2090 71 2490 118
rect 2090 37 2106 71
rect 2474 37 2490 71
rect 2090 21 2490 37
rect -2490 -37 -2090 -21
rect -2490 -71 -2474 -37
rect -2106 -71 -2090 -37
rect -2490 -118 -2090 -71
rect -2032 -37 -1632 -21
rect -2032 -71 -2016 -37
rect -1648 -71 -1632 -37
rect -2032 -118 -1632 -71
rect -1574 -37 -1174 -21
rect -1574 -71 -1558 -37
rect -1190 -71 -1174 -37
rect -1574 -118 -1174 -71
rect -1116 -37 -716 -21
rect -1116 -71 -1100 -37
rect -732 -71 -716 -37
rect -1116 -118 -716 -71
rect -658 -37 -258 -21
rect -658 -71 -642 -37
rect -274 -71 -258 -37
rect -658 -118 -258 -71
rect -200 -37 200 -21
rect -200 -71 -184 -37
rect 184 -71 200 -37
rect -200 -118 200 -71
rect 258 -37 658 -21
rect 258 -71 274 -37
rect 642 -71 658 -37
rect 258 -118 658 -71
rect 716 -37 1116 -21
rect 716 -71 732 -37
rect 1100 -71 1116 -37
rect 716 -118 1116 -71
rect 1174 -37 1574 -21
rect 1174 -71 1190 -37
rect 1558 -71 1574 -37
rect 1174 -118 1574 -71
rect 1632 -37 2032 -21
rect 1632 -71 1648 -37
rect 2016 -71 2032 -37
rect 1632 -118 2032 -71
rect 2090 -37 2490 -21
rect 2090 -71 2106 -37
rect 2474 -71 2490 -37
rect 2090 -118 2490 -71
rect -2490 -3365 -2090 -3318
rect -2490 -3399 -2474 -3365
rect -2106 -3399 -2090 -3365
rect -2490 -3415 -2090 -3399
rect -2032 -3365 -1632 -3318
rect -2032 -3399 -2016 -3365
rect -1648 -3399 -1632 -3365
rect -2032 -3415 -1632 -3399
rect -1574 -3365 -1174 -3318
rect -1574 -3399 -1558 -3365
rect -1190 -3399 -1174 -3365
rect -1574 -3415 -1174 -3399
rect -1116 -3365 -716 -3318
rect -1116 -3399 -1100 -3365
rect -732 -3399 -716 -3365
rect -1116 -3415 -716 -3399
rect -658 -3365 -258 -3318
rect -658 -3399 -642 -3365
rect -274 -3399 -258 -3365
rect -658 -3415 -258 -3399
rect -200 -3365 200 -3318
rect -200 -3399 -184 -3365
rect 184 -3399 200 -3365
rect -200 -3415 200 -3399
rect 258 -3365 658 -3318
rect 258 -3399 274 -3365
rect 642 -3399 658 -3365
rect 258 -3415 658 -3399
rect 716 -3365 1116 -3318
rect 716 -3399 732 -3365
rect 1100 -3399 1116 -3365
rect 716 -3415 1116 -3399
rect 1174 -3365 1574 -3318
rect 1174 -3399 1190 -3365
rect 1558 -3399 1574 -3365
rect 1174 -3415 1574 -3399
rect 1632 -3365 2032 -3318
rect 1632 -3399 1648 -3365
rect 2016 -3399 2032 -3365
rect 1632 -3415 2032 -3399
rect 2090 -3365 2490 -3318
rect 2090 -3399 2106 -3365
rect 2474 -3399 2490 -3365
rect 2090 -3415 2490 -3399
<< polycont >>
rect -2474 3365 -2106 3399
rect -2016 3365 -1648 3399
rect -1558 3365 -1190 3399
rect -1100 3365 -732 3399
rect -642 3365 -274 3399
rect -184 3365 184 3399
rect 274 3365 642 3399
rect 732 3365 1100 3399
rect 1190 3365 1558 3399
rect 1648 3365 2016 3399
rect 2106 3365 2474 3399
rect -2474 37 -2106 71
rect -2016 37 -1648 71
rect -1558 37 -1190 71
rect -1100 37 -732 71
rect -642 37 -274 71
rect -184 37 184 71
rect 274 37 642 71
rect 732 37 1100 71
rect 1190 37 1558 71
rect 1648 37 2016 71
rect 2106 37 2474 71
rect -2474 -71 -2106 -37
rect -2016 -71 -1648 -37
rect -1558 -71 -1190 -37
rect -1100 -71 -732 -37
rect -642 -71 -274 -37
rect -184 -71 184 -37
rect 274 -71 642 -37
rect 732 -71 1100 -37
rect 1190 -71 1558 -37
rect 1648 -71 2016 -37
rect 2106 -71 2474 -37
rect -2474 -3399 -2106 -3365
rect -2016 -3399 -1648 -3365
rect -1558 -3399 -1190 -3365
rect -1100 -3399 -732 -3365
rect -642 -3399 -274 -3365
rect -184 -3399 184 -3365
rect 274 -3399 642 -3365
rect 732 -3399 1100 -3365
rect 1190 -3399 1558 -3365
rect 1648 -3399 2016 -3365
rect 2106 -3399 2474 -3365
<< locali >>
rect -2650 3467 -2554 3501
rect 2554 3467 2650 3501
rect -2650 3405 -2616 3467
rect 2616 3405 2650 3467
rect -2490 3365 -2474 3399
rect -2106 3365 -2090 3399
rect -2032 3365 -2016 3399
rect -1648 3365 -1632 3399
rect -1574 3365 -1558 3399
rect -1190 3365 -1174 3399
rect -1116 3365 -1100 3399
rect -732 3365 -716 3399
rect -658 3365 -642 3399
rect -274 3365 -258 3399
rect -200 3365 -184 3399
rect 184 3365 200 3399
rect 258 3365 274 3399
rect 642 3365 658 3399
rect 716 3365 732 3399
rect 1100 3365 1116 3399
rect 1174 3365 1190 3399
rect 1558 3365 1574 3399
rect 1632 3365 1648 3399
rect 2016 3365 2032 3399
rect 2090 3365 2106 3399
rect 2474 3365 2490 3399
rect -2536 3306 -2502 3322
rect -2536 114 -2502 130
rect -2078 3306 -2044 3322
rect -2078 114 -2044 130
rect -1620 3306 -1586 3322
rect -1620 114 -1586 130
rect -1162 3306 -1128 3322
rect -1162 114 -1128 130
rect -704 3306 -670 3322
rect -704 114 -670 130
rect -246 3306 -212 3322
rect -246 114 -212 130
rect 212 3306 246 3322
rect 212 114 246 130
rect 670 3306 704 3322
rect 670 114 704 130
rect 1128 3306 1162 3322
rect 1128 114 1162 130
rect 1586 3306 1620 3322
rect 1586 114 1620 130
rect 2044 3306 2078 3322
rect 2044 114 2078 130
rect 2502 3306 2536 3322
rect 2502 114 2536 130
rect -2490 37 -2474 71
rect -2106 37 -2090 71
rect -2032 37 -2016 71
rect -1648 37 -1632 71
rect -1574 37 -1558 71
rect -1190 37 -1174 71
rect -1116 37 -1100 71
rect -732 37 -716 71
rect -658 37 -642 71
rect -274 37 -258 71
rect -200 37 -184 71
rect 184 37 200 71
rect 258 37 274 71
rect 642 37 658 71
rect 716 37 732 71
rect 1100 37 1116 71
rect 1174 37 1190 71
rect 1558 37 1574 71
rect 1632 37 1648 71
rect 2016 37 2032 71
rect 2090 37 2106 71
rect 2474 37 2490 71
rect -2490 -71 -2474 -37
rect -2106 -71 -2090 -37
rect -2032 -71 -2016 -37
rect -1648 -71 -1632 -37
rect -1574 -71 -1558 -37
rect -1190 -71 -1174 -37
rect -1116 -71 -1100 -37
rect -732 -71 -716 -37
rect -658 -71 -642 -37
rect -274 -71 -258 -37
rect -200 -71 -184 -37
rect 184 -71 200 -37
rect 258 -71 274 -37
rect 642 -71 658 -37
rect 716 -71 732 -37
rect 1100 -71 1116 -37
rect 1174 -71 1190 -37
rect 1558 -71 1574 -37
rect 1632 -71 1648 -37
rect 2016 -71 2032 -37
rect 2090 -71 2106 -37
rect 2474 -71 2490 -37
rect -2536 -130 -2502 -114
rect -2536 -3322 -2502 -3306
rect -2078 -130 -2044 -114
rect -2078 -3322 -2044 -3306
rect -1620 -130 -1586 -114
rect -1620 -3322 -1586 -3306
rect -1162 -130 -1128 -114
rect -1162 -3322 -1128 -3306
rect -704 -130 -670 -114
rect -704 -3322 -670 -3306
rect -246 -130 -212 -114
rect -246 -3322 -212 -3306
rect 212 -130 246 -114
rect 212 -3322 246 -3306
rect 670 -130 704 -114
rect 670 -3322 704 -3306
rect 1128 -130 1162 -114
rect 1128 -3322 1162 -3306
rect 1586 -130 1620 -114
rect 1586 -3322 1620 -3306
rect 2044 -130 2078 -114
rect 2044 -3322 2078 -3306
rect 2502 -130 2536 -114
rect 2502 -3322 2536 -3306
rect -2490 -3399 -2474 -3365
rect -2106 -3399 -2090 -3365
rect -2032 -3399 -2016 -3365
rect -1648 -3399 -1632 -3365
rect -1574 -3399 -1558 -3365
rect -1190 -3399 -1174 -3365
rect -1116 -3399 -1100 -3365
rect -732 -3399 -716 -3365
rect -658 -3399 -642 -3365
rect -274 -3399 -258 -3365
rect -200 -3399 -184 -3365
rect 184 -3399 200 -3365
rect 258 -3399 274 -3365
rect 642 -3399 658 -3365
rect 716 -3399 732 -3365
rect 1100 -3399 1116 -3365
rect 1174 -3399 1190 -3365
rect 1558 -3399 1574 -3365
rect 1632 -3399 1648 -3365
rect 2016 -3399 2032 -3365
rect 2090 -3399 2106 -3365
rect 2474 -3399 2490 -3365
rect -2650 -3467 -2616 -3405
rect 2616 -3467 2650 -3405
rect -2650 -3501 -2554 -3467
rect 2554 -3501 2650 -3467
<< viali >>
rect -2474 3365 -2106 3399
rect -2016 3365 -1648 3399
rect -1558 3365 -1190 3399
rect -1100 3365 -732 3399
rect -642 3365 -274 3399
rect -184 3365 184 3399
rect 274 3365 642 3399
rect 732 3365 1100 3399
rect 1190 3365 1558 3399
rect 1648 3365 2016 3399
rect 2106 3365 2474 3399
rect -2536 130 -2502 3306
rect -2078 130 -2044 3306
rect -1620 130 -1586 3306
rect -1162 130 -1128 3306
rect -704 130 -670 3306
rect -246 130 -212 3306
rect 212 130 246 3306
rect 670 130 704 3306
rect 1128 130 1162 3306
rect 1586 130 1620 3306
rect 2044 130 2078 3306
rect 2502 130 2536 3306
rect -2474 37 -2106 71
rect -2016 37 -1648 71
rect -1558 37 -1190 71
rect -1100 37 -732 71
rect -642 37 -274 71
rect -184 37 184 71
rect 274 37 642 71
rect 732 37 1100 71
rect 1190 37 1558 71
rect 1648 37 2016 71
rect 2106 37 2474 71
rect -2474 -71 -2106 -37
rect -2016 -71 -1648 -37
rect -1558 -71 -1190 -37
rect -1100 -71 -732 -37
rect -642 -71 -274 -37
rect -184 -71 184 -37
rect 274 -71 642 -37
rect 732 -71 1100 -37
rect 1190 -71 1558 -37
rect 1648 -71 2016 -37
rect 2106 -71 2474 -37
rect -2536 -3306 -2502 -130
rect -2078 -3306 -2044 -130
rect -1620 -3306 -1586 -130
rect -1162 -3306 -1128 -130
rect -704 -3306 -670 -130
rect -246 -3306 -212 -130
rect 212 -3306 246 -130
rect 670 -3306 704 -130
rect 1128 -3306 1162 -130
rect 1586 -3306 1620 -130
rect 2044 -3306 2078 -130
rect 2502 -3306 2536 -130
rect -2474 -3399 -2106 -3365
rect -2016 -3399 -1648 -3365
rect -1558 -3399 -1190 -3365
rect -1100 -3399 -732 -3365
rect -642 -3399 -274 -3365
rect -184 -3399 184 -3365
rect 274 -3399 642 -3365
rect 732 -3399 1100 -3365
rect 1190 -3399 1558 -3365
rect 1648 -3399 2016 -3365
rect 2106 -3399 2474 -3365
<< metal1 >>
rect -2486 3399 -2094 3405
rect -2486 3365 -2474 3399
rect -2106 3365 -2094 3399
rect -2486 3359 -2094 3365
rect -2028 3399 -1636 3405
rect -2028 3365 -2016 3399
rect -1648 3365 -1636 3399
rect -2028 3359 -1636 3365
rect -1570 3399 -1178 3405
rect -1570 3365 -1558 3399
rect -1190 3365 -1178 3399
rect -1570 3359 -1178 3365
rect -1112 3399 -720 3405
rect -1112 3365 -1100 3399
rect -732 3365 -720 3399
rect -1112 3359 -720 3365
rect -654 3399 -262 3405
rect -654 3365 -642 3399
rect -274 3365 -262 3399
rect -654 3359 -262 3365
rect -196 3399 196 3405
rect -196 3365 -184 3399
rect 184 3365 196 3399
rect -196 3359 196 3365
rect 262 3399 654 3405
rect 262 3365 274 3399
rect 642 3365 654 3399
rect 262 3359 654 3365
rect 720 3399 1112 3405
rect 720 3365 732 3399
rect 1100 3365 1112 3399
rect 720 3359 1112 3365
rect 1178 3399 1570 3405
rect 1178 3365 1190 3399
rect 1558 3365 1570 3399
rect 1178 3359 1570 3365
rect 1636 3399 2028 3405
rect 1636 3365 1648 3399
rect 2016 3365 2028 3399
rect 1636 3359 2028 3365
rect 2094 3399 2486 3405
rect 2094 3365 2106 3399
rect 2474 3365 2486 3399
rect 2094 3359 2486 3365
rect -2542 3306 -2496 3318
rect -2542 130 -2536 3306
rect -2502 130 -2496 3306
rect -2542 118 -2496 130
rect -2084 3306 -2038 3318
rect -2084 130 -2078 3306
rect -2044 130 -2038 3306
rect -2084 118 -2038 130
rect -1626 3306 -1580 3318
rect -1626 130 -1620 3306
rect -1586 130 -1580 3306
rect -1626 118 -1580 130
rect -1168 3306 -1122 3318
rect -1168 130 -1162 3306
rect -1128 130 -1122 3306
rect -1168 118 -1122 130
rect -710 3306 -664 3318
rect -710 130 -704 3306
rect -670 130 -664 3306
rect -710 118 -664 130
rect -252 3306 -206 3318
rect -252 130 -246 3306
rect -212 130 -206 3306
rect -252 118 -206 130
rect 206 3306 252 3318
rect 206 130 212 3306
rect 246 130 252 3306
rect 206 118 252 130
rect 664 3306 710 3318
rect 664 130 670 3306
rect 704 130 710 3306
rect 664 118 710 130
rect 1122 3306 1168 3318
rect 1122 130 1128 3306
rect 1162 130 1168 3306
rect 1122 118 1168 130
rect 1580 3306 1626 3318
rect 1580 130 1586 3306
rect 1620 130 1626 3306
rect 1580 118 1626 130
rect 2038 3306 2084 3318
rect 2038 130 2044 3306
rect 2078 130 2084 3306
rect 2038 118 2084 130
rect 2496 3306 2542 3318
rect 2496 130 2502 3306
rect 2536 130 2542 3306
rect 2496 118 2542 130
rect -2486 71 -2094 77
rect -2486 37 -2474 71
rect -2106 37 -2094 71
rect -2486 31 -2094 37
rect -2028 71 -1636 77
rect -2028 37 -2016 71
rect -1648 37 -1636 71
rect -2028 31 -1636 37
rect -1570 71 -1178 77
rect -1570 37 -1558 71
rect -1190 37 -1178 71
rect -1570 31 -1178 37
rect -1112 71 -720 77
rect -1112 37 -1100 71
rect -732 37 -720 71
rect -1112 31 -720 37
rect -654 71 -262 77
rect -654 37 -642 71
rect -274 37 -262 71
rect -654 31 -262 37
rect -196 71 196 77
rect -196 37 -184 71
rect 184 37 196 71
rect -196 31 196 37
rect 262 71 654 77
rect 262 37 274 71
rect 642 37 654 71
rect 262 31 654 37
rect 720 71 1112 77
rect 720 37 732 71
rect 1100 37 1112 71
rect 720 31 1112 37
rect 1178 71 1570 77
rect 1178 37 1190 71
rect 1558 37 1570 71
rect 1178 31 1570 37
rect 1636 71 2028 77
rect 1636 37 1648 71
rect 2016 37 2028 71
rect 1636 31 2028 37
rect 2094 71 2486 77
rect 2094 37 2106 71
rect 2474 37 2486 71
rect 2094 31 2486 37
rect -2486 -37 -2094 -31
rect -2486 -71 -2474 -37
rect -2106 -71 -2094 -37
rect -2486 -77 -2094 -71
rect -2028 -37 -1636 -31
rect -2028 -71 -2016 -37
rect -1648 -71 -1636 -37
rect -2028 -77 -1636 -71
rect -1570 -37 -1178 -31
rect -1570 -71 -1558 -37
rect -1190 -71 -1178 -37
rect -1570 -77 -1178 -71
rect -1112 -37 -720 -31
rect -1112 -71 -1100 -37
rect -732 -71 -720 -37
rect -1112 -77 -720 -71
rect -654 -37 -262 -31
rect -654 -71 -642 -37
rect -274 -71 -262 -37
rect -654 -77 -262 -71
rect -196 -37 196 -31
rect -196 -71 -184 -37
rect 184 -71 196 -37
rect -196 -77 196 -71
rect 262 -37 654 -31
rect 262 -71 274 -37
rect 642 -71 654 -37
rect 262 -77 654 -71
rect 720 -37 1112 -31
rect 720 -71 732 -37
rect 1100 -71 1112 -37
rect 720 -77 1112 -71
rect 1178 -37 1570 -31
rect 1178 -71 1190 -37
rect 1558 -71 1570 -37
rect 1178 -77 1570 -71
rect 1636 -37 2028 -31
rect 1636 -71 1648 -37
rect 2016 -71 2028 -37
rect 1636 -77 2028 -71
rect 2094 -37 2486 -31
rect 2094 -71 2106 -37
rect 2474 -71 2486 -37
rect 2094 -77 2486 -71
rect -2542 -130 -2496 -118
rect -2542 -3306 -2536 -130
rect -2502 -3306 -2496 -130
rect -2542 -3318 -2496 -3306
rect -2084 -130 -2038 -118
rect -2084 -3306 -2078 -130
rect -2044 -3306 -2038 -130
rect -2084 -3318 -2038 -3306
rect -1626 -130 -1580 -118
rect -1626 -3306 -1620 -130
rect -1586 -3306 -1580 -130
rect -1626 -3318 -1580 -3306
rect -1168 -130 -1122 -118
rect -1168 -3306 -1162 -130
rect -1128 -3306 -1122 -130
rect -1168 -3318 -1122 -3306
rect -710 -130 -664 -118
rect -710 -3306 -704 -130
rect -670 -3306 -664 -130
rect -710 -3318 -664 -3306
rect -252 -130 -206 -118
rect -252 -3306 -246 -130
rect -212 -3306 -206 -130
rect -252 -3318 -206 -3306
rect 206 -130 252 -118
rect 206 -3306 212 -130
rect 246 -3306 252 -130
rect 206 -3318 252 -3306
rect 664 -130 710 -118
rect 664 -3306 670 -130
rect 704 -3306 710 -130
rect 664 -3318 710 -3306
rect 1122 -130 1168 -118
rect 1122 -3306 1128 -130
rect 1162 -3306 1168 -130
rect 1122 -3318 1168 -3306
rect 1580 -130 1626 -118
rect 1580 -3306 1586 -130
rect 1620 -3306 1626 -130
rect 1580 -3318 1626 -3306
rect 2038 -130 2084 -118
rect 2038 -3306 2044 -130
rect 2078 -3306 2084 -130
rect 2038 -3318 2084 -3306
rect 2496 -130 2542 -118
rect 2496 -3306 2502 -130
rect 2536 -3306 2542 -130
rect 2496 -3318 2542 -3306
rect -2486 -3365 -2094 -3359
rect -2486 -3399 -2474 -3365
rect -2106 -3399 -2094 -3365
rect -2486 -3405 -2094 -3399
rect -2028 -3365 -1636 -3359
rect -2028 -3399 -2016 -3365
rect -1648 -3399 -1636 -3365
rect -2028 -3405 -1636 -3399
rect -1570 -3365 -1178 -3359
rect -1570 -3399 -1558 -3365
rect -1190 -3399 -1178 -3365
rect -1570 -3405 -1178 -3399
rect -1112 -3365 -720 -3359
rect -1112 -3399 -1100 -3365
rect -732 -3399 -720 -3365
rect -1112 -3405 -720 -3399
rect -654 -3365 -262 -3359
rect -654 -3399 -642 -3365
rect -274 -3399 -262 -3365
rect -654 -3405 -262 -3399
rect -196 -3365 196 -3359
rect -196 -3399 -184 -3365
rect 184 -3399 196 -3365
rect -196 -3405 196 -3399
rect 262 -3365 654 -3359
rect 262 -3399 274 -3365
rect 642 -3399 654 -3365
rect 262 -3405 654 -3399
rect 720 -3365 1112 -3359
rect 720 -3399 732 -3365
rect 1100 -3399 1112 -3365
rect 720 -3405 1112 -3399
rect 1178 -3365 1570 -3359
rect 1178 -3399 1190 -3365
rect 1558 -3399 1570 -3365
rect 1178 -3405 1570 -3399
rect 1636 -3365 2028 -3359
rect 1636 -3399 1648 -3365
rect 2016 -3399 2028 -3365
rect 1636 -3405 2028 -3399
rect 2094 -3365 2486 -3359
rect 2094 -3399 2106 -3365
rect 2474 -3399 2486 -3365
rect 2094 -3405 2486 -3399
<< properties >>
string FIXED_BBOX -2633 -3484 2633 3484
string gencell sky130_fd_pr__pfet_01v8_lvt
string library sky130
string parameters w 16 l 2 m 2 nf 11 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.35 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
