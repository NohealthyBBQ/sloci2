magic
tech sky130A
magscale 1 2
timestamp 1672354881
<< locali >>
rect 3500 -3700 4020 -3000
rect 3500 -4200 3800 -3700
rect 4000 -4200 4020 -3700
rect 3500 -4980 4020 -4200
rect 12280 -60200 12320 -60140
rect 17840 -60160 23140 -60120
rect 12280 -60260 13060 -60200
rect 17840 -60260 17940 -60160
rect 18920 -60260 22060 -60160
rect 23040 -60260 23140 -60160
rect 17840 -60300 23140 -60260
<< viali >>
rect 3800 -4200 4000 -3700
rect 17940 -60260 18920 -60160
rect 22060 -60260 23040 -60160
<< metal1 >>
rect -960 3080 60 3100
rect -960 2980 -940 3080
rect -840 2980 60 3080
rect -960 2960 60 2980
rect 890 2660 900 2860
rect 1100 2660 1110 2860
rect -60 2160 100 2180
rect -60 2060 -40 2160
rect 60 2060 100 2160
rect -60 2040 100 2060
rect -300 1860 300 1900
rect -300 1740 -260 1860
rect -140 1740 300 1860
rect -300 1700 300 1740
rect 260 1380 540 1480
rect 260 1280 280 1380
rect 520 1280 540 1380
rect 260 1260 540 1280
rect 3380 -2380 3560 -2360
rect 3380 -2440 3480 -2380
rect 3540 -2440 3560 -2380
rect 3380 -2460 3560 -2440
rect 3794 -3700 4006 -3688
rect 3790 -4200 3800 -3700
rect 4000 -4200 4010 -3700
rect 3794 -4212 4006 -4200
rect 3260 -5220 3420 -4560
rect 3260 -5340 3280 -5220
rect 3400 -5340 3420 -5220
rect 3260 -5380 3420 -5340
rect -960 -24920 360 -24900
rect -960 -25020 -940 -24920
rect -840 -25020 360 -24920
rect -960 -25040 360 -25020
rect 1070 -25320 1080 -25120
rect 1360 -25320 1370 -25120
rect -580 -25840 300 -25820
rect -580 -25940 -560 -25840
rect -420 -25940 300 -25840
rect -580 -25960 300 -25940
rect -340 -26160 520 -26120
rect -340 -26340 -300 -26160
rect -160 -26340 520 -26160
rect -340 -26380 520 -26340
rect -960 -52520 220 -52500
rect -960 -52620 -940 -52520
rect -840 -52620 220 -52520
rect -960 -52640 220 -52620
rect 990 -53000 1000 -52800
rect 1200 -53000 1210 -52800
rect -60 -53440 80 -53420
rect -60 -53540 -40 -53440
rect 60 -53540 80 -53440
rect -60 -53560 80 -53540
rect -340 -53780 320 -53740
rect -340 -53940 -300 -53780
rect -160 -53940 320 -53780
rect -340 -53980 320 -53940
rect 11820 -54640 12280 -54630
rect 11820 -54700 12180 -54640
rect 12260 -54700 12280 -54640
rect 11820 -54710 12280 -54700
rect 12160 -58460 12780 -58440
rect 12160 -58600 12180 -58460
rect 12260 -58600 12780 -58460
rect 12160 -58620 12780 -58600
rect 12870 -59340 12880 -59140
rect 12940 -59340 12950 -59140
rect 17928 -60160 18932 -60154
rect 17928 -60260 17940 -60160
rect 18920 -60260 18932 -60160
rect 17928 -60266 18932 -60260
rect 22048 -60160 23052 -60154
rect 22048 -60260 22060 -60160
rect 23040 -60260 23052 -60160
rect 22048 -60266 23052 -60260
<< via1 >>
rect -940 2980 -840 3080
rect 900 2660 1100 2860
rect -40 2060 60 2160
rect -260 1740 -140 1860
rect 280 1280 520 1380
rect 3480 -2440 3540 -2380
rect 3800 -4200 4000 -3700
rect 3280 -5340 3400 -5220
rect -940 -25020 -840 -24920
rect 1080 -25320 1360 -25120
rect -560 -25940 -420 -25840
rect -300 -26340 -160 -26160
rect -940 -52620 -840 -52520
rect 1000 -53000 1200 -52800
rect -40 -53540 60 -53440
rect -300 -53940 -160 -53780
rect 12180 -54700 12260 -54640
rect 12180 -58600 12260 -58460
rect 12880 -59340 12940 -59140
rect 17940 -60260 18920 -60160
rect 22060 -60260 23040 -60160
<< metal2 >>
rect -1100 3080 -700 3200
rect -1100 2980 -940 3080
rect -840 2980 -700 3080
rect -1100 -24920 -700 2980
rect 900 2860 1100 2870
rect 900 2650 1100 2660
rect -60 2160 80 2180
rect -60 2060 -40 2160
rect 60 2060 80 2160
rect -260 1860 -140 1870
rect -260 1730 -140 1740
rect -60 -1000 80 2060
rect 280 1380 520 1390
rect 280 1270 520 1280
rect -60 -1140 3560 -1000
rect 3460 -2380 3560 -1140
rect 3460 -2440 3480 -2380
rect 3540 -2440 3560 -2380
rect 3460 -2460 3560 -2440
rect 3340 -3440 3680 -3280
rect 3540 -5000 3680 -3440
rect 3800 -3700 4000 -3690
rect 3800 -4210 4000 -4200
rect -1100 -25020 -940 -24920
rect -840 -25020 -700 -24920
rect -1100 -52520 -700 -25020
rect -560 -5140 3680 -5000
rect -560 -25840 -420 -5140
rect -560 -25960 -420 -25940
rect -60 -5220 3420 -5200
rect -60 -5340 3280 -5220
rect 3400 -5340 3420 -5220
rect -60 -5360 3420 -5340
rect -300 -26160 -160 -26150
rect -300 -26350 -160 -26340
rect -1100 -52620 -940 -52520
rect -840 -52620 -700 -52520
rect -1100 -52700 -700 -52620
rect -60 -53440 80 -5360
rect 1080 -25120 1360 -25110
rect 1080 -25330 1360 -25320
rect 1000 -52800 1200 -52790
rect 1000 -53010 1200 -53000
rect 10200 -53000 10600 -52900
rect -60 -53540 -40 -53440
rect 60 -53540 80 -53440
rect -60 -53560 80 -53540
rect 10200 -53500 10300 -53000
rect 10500 -53500 10600 -53000
rect 10200 -53600 10600 -53500
rect 19200 -53200 19500 -53190
rect 19200 -53510 19500 -53500
rect -300 -53780 -160 -53760
rect -300 -57080 -160 -53940
rect 12180 -54640 12260 -54630
rect -300 -57100 3040 -57080
rect -300 -57180 2940 -57100
rect 3020 -57180 3040 -57100
rect -300 -57200 3040 -57180
rect 12180 -58460 12260 -54700
rect 2880 -58560 3020 -58540
rect 2880 -58640 2940 -58560
rect 12180 -58620 12260 -58600
rect 2880 -58660 3020 -58640
rect 2880 -58760 3020 -58740
rect 2880 -58840 2940 -58760
rect 2880 -58860 3020 -58840
rect 3400 -58760 4160 -58700
rect 3480 -58860 4160 -58760
rect 3400 -58880 4160 -58860
rect 6300 -59140 12960 -59100
rect 6300 -59340 12880 -59140
rect 12940 -59340 12960 -59140
rect 6300 -59400 12960 -59340
rect 17940 -60160 18920 -60150
rect 17940 -60270 18920 -60260
rect 22060 -60160 23040 -60150
rect 22060 -60270 23040 -60260
<< via2 >>
rect 900 2660 1100 2860
rect -260 1740 -140 1860
rect 280 1280 520 1380
rect 3800 -4200 4000 -3700
rect -300 -26340 -160 -26160
rect 1080 -25320 1360 -25120
rect 1000 -53000 1200 -52800
rect 10300 -53500 10500 -53000
rect 19200 -53500 19500 -53200
rect -300 -53940 -160 -53780
rect 2940 -57180 3020 -57100
rect 2940 -58640 3020 -58560
rect 2940 -58840 3020 -58760
rect 3400 -58860 3480 -58760
rect 17940 -60260 18920 -60160
rect 22060 -60260 23040 -60160
<< metal3 >>
rect 890 2860 1110 2865
rect 890 2660 900 2860
rect 1100 2660 1110 2860
rect 890 2655 1110 2660
rect -380 1860 -100 2440
rect -380 1740 -260 1860
rect -140 1740 -100 1860
rect -380 -26160 -100 1740
rect 200 1380 600 1400
rect 200 1280 280 1380
rect 520 1280 600 1380
rect 200 -200 600 1280
rect 200 -800 7000 -200
rect 3780 -3700 6780 -3680
rect 3780 -4200 3800 -3700
rect 4000 -4200 6780 -3700
rect 3780 -4220 6780 -4200
rect 1070 -25120 1370 -25115
rect 1070 -25320 1080 -25120
rect 1360 -25320 1370 -25120
rect 1070 -25325 1370 -25320
rect -380 -26340 -300 -26160
rect -160 -26340 -100 -26160
rect -380 -53100 -100 -26340
rect 990 -52800 1210 -52795
rect 990 -53000 1000 -52800
rect 1200 -53000 1210 -52800
rect 990 -53005 1210 -53000
rect 10290 -53000 10510 -52995
rect 4060 -53100 4420 -53060
rect 10290 -53100 10300 -53000
rect -380 -53400 4420 -53100
rect -380 -53780 -100 -53400
rect 4060 -53680 4420 -53400
rect 10200 -53500 10300 -53100
rect 10500 -53100 10510 -53000
rect 10500 -53200 19600 -53100
rect 10500 -53500 19200 -53200
rect 19500 -53500 19600 -53200
rect 10200 -53600 19600 -53500
rect -380 -53940 -300 -53780
rect -160 -53940 -100 -53780
rect -380 -54040 -100 -53940
rect 2920 -57100 3040 -57080
rect 2920 -57180 2940 -57100
rect 3020 -57180 3040 -57100
rect 2920 -58560 3040 -57180
rect 2920 -58640 2940 -58560
rect 3020 -58640 3040 -58560
rect 2920 -58660 3040 -58640
rect 2920 -58760 3500 -58740
rect 2920 -58840 2940 -58760
rect 3020 -58840 3400 -58760
rect 2920 -58860 3400 -58840
rect 3480 -58860 3500 -58760
rect 2920 -58880 3500 -58860
rect 17910 -60300 17920 -60140
rect 18940 -60300 18950 -60140
rect 22030 -60280 22040 -60140
rect 23060 -60280 23070 -60140
<< via3 >>
rect 900 2660 1100 2860
rect 1080 -25320 1360 -25120
rect 1000 -53000 1200 -52800
rect 17920 -60160 18940 -60140
rect 17920 -60260 17940 -60160
rect 17940 -60260 18920 -60160
rect 18920 -60260 18940 -60160
rect 17920 -60300 18940 -60260
rect 22040 -60160 23060 -60140
rect 22040 -60260 22060 -60160
rect 22060 -60260 23040 -60160
rect 23040 -60260 23060 -60160
rect 22040 -60280 23060 -60260
<< metal4 >>
rect 6200 27400 25600 28600
rect 800 3000 5400 3200
rect 800 2860 1200 3000
rect 800 2660 900 2860
rect 1100 2660 1200 2860
rect 800 2600 1200 2660
rect 24800 -4600 25600 27400
rect 12800 -5400 25600 -4600
rect 1020 -25000 5340 -24800
rect 1020 -25120 1440 -25000
rect 1020 -25320 1080 -25120
rect 1360 -25320 1440 -25120
rect 1020 -25360 1440 -25320
rect 24800 -32200 25600 -5400
rect 12800 -33000 25600 -32200
rect 1000 -52600 5200 -52400
rect 1000 -52799 1200 -52600
rect 999 -52800 1201 -52799
rect 999 -53000 1000 -52800
rect 1200 -53000 1201 -52800
rect 999 -53001 1201 -53000
rect 200 -60600 12320 -60200
rect 17380 -60600 17520 -59780
rect 17840 -60140 23140 -60120
rect 17840 -60300 17920 -60140
rect 18940 -60280 22040 -60140
rect 23060 -60200 23140 -60140
rect 24800 -60200 25600 -33000
rect 23060 -60280 25600 -60200
rect 18940 -60300 25600 -60280
rect 17840 -60600 25600 -60300
rect 200 -61000 25600 -60600
use 2_to_4_decoder  2_to_4_decoder_0
timestamp 1671728743
transform 1 0 1060 0 1 -3080
box -460 -1920 2480 1848
use 3T  3T_0
timestamp 1671680485
transform 1 0 280 0 1 2300
box -280 -900 1153 838
use 3T  3T_1
timestamp 1671680485
transform 1 0 280 0 1 -53300
box -280 -900 1153 838
use 3T  3T_2
timestamp 1671680485
transform 1 0 480 0 1 -25700
box -280 -900 1153 838
use bias  bias_0
timestamp 1672278816
transform 1 0 17763 0 1 -60200
box 37 -200 5412 8450
use cd_current  cd_current_0
timestamp 1672331172
transform 1 0 1300 0 1 -54260
box 40 -200 5412 1200
use cd_output  cd_output_0
timestamp 1672344752
transform 1 0 8673 0 1 -54767
box -53 -53 3441 1915
use opamp_realcomp3_usefinger  opamp_realcomp3_usefinger_0
timestamp 1662739988
transform 1 0 5580 0 1 -60994
box -5380 594 6776 6403
use rc_model_4cap  rc_model_4cap_0
timestamp 1672330275
transform 1 0 -8000 0 1 19400
box 8000 -16400 25896 9200
use rc_model_6cap  rc_model_6cap_0
timestamp 1672329859
transform 1 0 -1400 0 1 -8600
box 1400 -16400 25896 9200
use rc_model_8cap  rc_model_8cap_0
timestamp 1672329920
transform 1 0 -1406 0 1 -36198
box 1400 -16400 25896 9200
use sample_hold  sample_hold_0
timestamp 1672262444
transform 1 0 7400 0 1 -60200
box 5200 -200 10099 4000
<< labels >>
flabel metal4 800 2860 1200 3200 0 FreeSans 1600 0 0 0 Vin_1
flabel metal4 1020 -25120 1440 -24800 0 FreeSans 1600 0 0 0 Vin_2
flabel metal4 1000 -52800 1200 -52400 0 FreeSans 1600 0 0 0 Vin_3
flabel metal2 -60 -1140 3560 -1000 0 FreeSans 1600 0 0 0 D1
flabel metal2 -560 -5140 3680 -5000 0 FreeSans 1600 0 0 0 D2
flabel metal2 -60 -5360 3280 -5200 0 FreeSans 1600 0 0 0 D3
flabel metal3 -380 -53780 -100 -26340 0 FreeSans 1600 0 0 0 Vpixel_out
flabel space 6204 -59400 12880 -59100 0 FreeSans 1600 0 0 0 Vbuff_out
<< end >>
