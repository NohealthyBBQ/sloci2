magic
tech sky130A
magscale 1 2
timestamp 1662836520
<< locali >>
rect -5320 3700 -2040 3760
rect -5320 3600 -5220 3700
rect -5320 3200 -5300 3600
rect -5240 3200 -5220 3600
rect -5320 2500 -5220 3200
rect -5320 2100 -5300 2500
rect -5240 2100 -5220 2500
rect -5320 1380 -5220 2100
rect -5320 980 -5300 1380
rect -5240 980 -5220 1380
rect -5320 820 -5220 980
rect -4080 900 -4000 3700
rect -4080 820 -2040 900
<< viali >>
rect -5300 3200 -5240 3600
rect -5300 2100 -5240 2500
rect -5300 980 -5240 1380
rect 4820 780 5140 860
<< metal1 >>
rect -5170 5620 -5160 5680
rect -4760 5620 -4750 5680
rect -3730 5620 -3720 5680
rect -3320 5620 -3310 5680
rect -2690 5620 -2680 5680
rect -2280 5620 -2270 5680
rect -1230 5620 -1220 5680
rect -820 5620 -810 5680
rect -5170 4040 -5160 4100
rect -4760 4040 -4750 4100
rect -3730 4044 -3720 4100
rect -3320 4044 -3310 4100
rect -2272 4044 -2270 4100
rect -1230 4040 -1220 4100
rect -820 4040 -810 4100
rect -5306 3600 -5234 3612
rect -5310 3200 -5300 3600
rect -5240 3200 -5230 3600
rect -4100 3240 -3980 3720
rect -5306 3188 -5234 3200
rect -4100 2840 -4060 3240
rect -4000 2840 -3980 3240
rect -5306 2500 -5234 2512
rect -5310 2100 -5300 2500
rect -5240 2100 -5230 2500
rect -4100 2120 -3980 2840
rect 510 2600 520 2660
rect 580 2600 590 2660
rect -5306 2088 -5234 2100
rect -4100 1720 -4060 2120
rect -4000 1720 -3980 2120
rect -5306 1380 -5234 1392
rect -5310 980 -5300 1380
rect -5240 980 -5230 1380
rect -5306 968 -5234 980
rect -4685 770 -4625 966
rect -4100 880 -3980 1720
rect 6290 1100 6300 1400
rect 6500 1100 6510 1400
rect 3346 966 3356 1031
rect -3470 880 -3460 940
rect -2760 880 -2750 940
rect 3338 928 3356 966
rect 3431 963 3441 1031
rect 3431 928 3459 963
rect 3338 907 3459 928
rect 4808 860 5152 866
rect 4808 780 4820 860
rect 5140 780 5152 860
rect 4808 774 5152 780
rect -4685 710 -750 770
rect -4685 701 -4625 710
rect -1324 594 -1276 710
<< via1 >>
rect -5160 5620 -4760 5680
rect -3720 5620 -3320 5680
rect -2680 5620 -2280 5680
rect -1220 5620 -820 5680
rect -5160 4040 -4760 4100
rect -1220 4040 -820 4100
rect -5300 3200 -5240 3600
rect -4060 2840 -4000 3240
rect -5300 2100 -5240 2500
rect 520 2600 580 2660
rect -4060 1720 -4000 2120
rect -5300 980 -5240 1380
rect 6300 1100 6500 1400
rect -3460 880 -2760 940
rect 3356 928 3431 1031
rect 4820 780 5140 860
<< metal2 >>
rect -5160 5680 -4760 5690
rect -5160 5610 -4760 5620
rect -3720 5680 -3320 5690
rect -3720 5610 -3320 5620
rect -2680 5680 -2280 5690
rect -2680 5610 -2280 5620
rect -1220 5680 -820 5690
rect -1220 5610 -820 5620
rect -5160 4100 -4760 4110
rect -5160 4030 -4760 4040
rect -1220 4100 -820 4110
rect -1220 4030 -820 4040
rect 300 3670 650 3800
rect -5300 3600 -5240 3610
rect -5300 3190 -5240 3200
rect -4060 3240 -4000 3250
rect 280 2913 736 3045
rect -4060 2830 -4000 2840
rect -3780 2660 -3710 2670
rect -3780 2590 -3710 2600
rect -2480 2660 590 2670
rect -2480 2600 -1740 2660
rect -1670 2600 520 2660
rect 580 2600 590 2660
rect -2480 2590 590 2600
rect -5300 2500 -5240 2510
rect -2752 2352 -2652 2432
rect -4080 2330 -4000 2340
rect -4080 2260 -4000 2270
rect -2752 2172 -2652 2252
rect 301 2157 647 2289
rect -5300 2090 -5240 2100
rect -4060 2120 -4000 2130
rect -4060 1710 -4000 1720
rect 305 1401 651 1533
rect 6300 1400 6500 1410
rect -5300 1380 -5240 1390
rect 6300 1090 6500 1100
rect -5300 970 -5240 980
rect 3009 1031 3459 1047
rect -3460 940 -2760 950
rect 3009 928 3356 1031
rect 3431 928 3459 1031
rect 3009 907 3459 928
rect -3460 800 -2760 880
rect 4820 860 5140 870
rect 4820 770 5140 780
rect -3460 730 -2760 740
<< via2 >>
rect -5160 5620 -4760 5680
rect -3720 5620 -3320 5680
rect -2680 5620 -2280 5680
rect -1220 5620 -820 5680
rect -5160 4040 -4760 4100
rect -1220 4040 -820 4100
rect -5300 3200 -5240 3600
rect -4060 2840 -4000 3240
rect -3780 2600 -3710 2660
rect -1740 2600 -1670 2660
rect -5300 2100 -5240 2500
rect -4080 2270 -4000 2330
rect -4060 1720 -4000 2120
rect -5300 980 -5240 1380
rect 6300 1100 6500 1400
rect -3460 740 -2760 800
rect 4820 780 5140 860
<< metal3 >>
rect -5170 5620 -5160 5720
rect -4760 5620 -4750 5720
rect -5170 5615 -4750 5620
rect -3730 5620 -3720 5720
rect -3320 5620 -3310 5720
rect -3730 5615 -3310 5620
rect -2690 5620 -2680 5720
rect -2280 5620 -2270 5720
rect -2690 5615 -2270 5620
rect -1230 5620 -1220 5720
rect -820 5620 -810 5720
rect 1810 5620 1820 5780
rect 1940 5620 1950 5780
rect -1230 5615 -810 5620
rect -1750 4874 -1740 4950
rect -1664 4874 -1654 4950
rect -5170 4100 -4750 4105
rect -5170 4000 -5160 4100
rect -4760 4000 -4750 4100
rect -5310 3600 -5230 3605
rect -5350 3200 -5340 3600
rect -5240 3200 -5230 3600
rect -5310 3195 -5230 3200
rect -4070 3240 -3990 3245
rect -4070 2840 -4060 3240
rect -3960 2840 -3950 3240
rect -4070 2835 -3990 2840
rect -3832 2660 -3700 4300
rect -1230 4100 -810 4105
rect -3832 2600 -3780 2660
rect -3710 2600 -3700 2660
rect -3832 2590 -3700 2600
rect -1772 2660 -1642 4038
rect -1230 4000 -1220 4100
rect -820 4000 -810 4100
rect 1810 3920 1820 4100
rect 1940 3920 1950 4100
rect -1772 2600 -1740 2660
rect -1670 2600 -1642 2660
rect -1772 2560 -1642 2600
rect -5310 2500 -5230 2505
rect -5350 2100 -5340 2500
rect -5240 2100 -5230 2500
rect -4090 2330 -3990 2335
rect -4090 2270 -4080 2330
rect -4000 2270 -3990 2330
rect -4090 2265 -3990 2270
rect -5310 2095 -5230 2100
rect -4070 2120 -3990 2125
rect -4070 1720 -4060 2120
rect -3960 1720 -3950 2120
rect -4070 1715 -3990 1720
rect 6300 1405 6500 1800
rect 6290 1400 6510 1405
rect -5310 1380 -5230 1385
rect -5350 980 -5340 1380
rect -5240 980 -5230 1380
rect 6290 1100 6300 1400
rect 6500 1100 6510 1400
rect 6290 1095 6510 1100
rect -5310 975 -5230 980
rect 4810 860 5150 865
rect -3470 740 -3460 840
rect -2760 740 -2750 840
rect -3470 735 -2750 740
rect -1080 720 -1070 850
rect -970 720 -960 850
rect 4810 740 4820 860
rect 5140 740 5150 860
<< via3 >>
rect -5160 5680 -4760 5720
rect -5160 5620 -4760 5680
rect -3720 5680 -3320 5720
rect -3720 5620 -3320 5680
rect -2680 5680 -2280 5720
rect -2680 5620 -2280 5680
rect -1220 5680 -820 5720
rect -1220 5620 -820 5680
rect 1820 5620 1940 5780
rect -1740 4874 -1664 4950
rect -5160 4040 -4760 4100
rect -5160 4000 -4760 4040
rect -5340 3200 -5300 3600
rect -5300 3200 -5240 3600
rect -4060 2840 -4000 3240
rect -4000 2840 -3960 3240
rect -1220 4040 -820 4100
rect -1220 4000 -820 4040
rect 1820 3940 1940 4100
rect -5340 2100 -5300 2500
rect -5300 2100 -5240 2500
rect -4060 1720 -4000 2120
rect -4000 1720 -3960 2120
rect -5340 980 -5300 1380
rect -5300 980 -5240 1380
rect -3460 800 -2760 840
rect -3460 740 -2760 800
rect -1070 720 -970 850
rect 4820 780 5140 860
rect 4820 740 5140 780
<< metal4 >>
rect -5380 5780 3000 5800
rect -5380 5720 1820 5780
rect -5380 5620 -5160 5720
rect -4760 5620 -3720 5720
rect -3320 5620 -2680 5720
rect -2280 5620 -1220 5720
rect -820 5620 1820 5720
rect 1940 5620 3000 5780
rect -5380 5600 3000 5620
rect -5380 4120 -5180 5600
rect -1741 4950 -1663 4951
rect -1741 4874 -1740 4950
rect -1664 4940 -1663 4950
rect -1664 4880 3520 4940
rect -1664 4874 -1663 4880
rect -1741 4873 -1663 4874
rect -5380 4100 3000 4120
rect -5380 4000 -5160 4100
rect -4760 4000 -1220 4100
rect -820 4000 1820 4100
rect -5380 3940 1820 4000
rect 1940 3940 3000 4100
rect -5380 3920 3000 3940
rect -5380 3600 3160 3800
rect -5380 3200 -5340 3600
rect -5240 3200 -5180 3600
rect -5380 2500 -5180 3200
rect -5380 2100 -5340 2500
rect -5240 2100 -5180 2500
rect -5380 1380 -5180 2100
rect -5380 980 -5340 1380
rect -5240 980 -5180 1380
rect -5380 860 -5180 980
rect -4100 3240 -3900 3600
rect -4100 2840 -4060 3240
rect -3960 2840 -3900 3240
rect -4100 2120 -3900 2840
rect -4100 1720 -4060 2120
rect -3960 1720 -3900 2120
rect -4100 860 -3900 1720
rect 4819 860 5141 861
rect -5380 850 4820 860
rect -5380 840 -1070 850
rect -5380 740 -3460 840
rect -2760 740 -1070 840
rect -5380 720 -1070 740
rect -970 740 4820 850
rect 5140 740 6740 860
rect -970 720 6740 740
rect -5380 660 6740 720
use XM_actload2  XM_actload2_0
timestamp 1662836520
transform 1 0 -2047 0 1 753
box -53 -53 2571 3173
use XM_cs  XM_cs_0
timestamp 1662401230
transform 1 0 664 0 1 753
box -140 -53 2482 5650
use XM_diffpair  XM_diffpair_0
timestamp 1662590620
transform 1 0 -3688 0 1 2162
box -400 -1400 1600 1700
use XM_ppair  XM_ppair_0
timestamp 1662597113
transform 1 0 -5102 0 1 5030
box -220 -1060 4440 720
use XM_tail  XM_tail_0
timestamp 1662390953
transform 1 0 -5225 0 1 839
box -53 -51 1200 2931
use sky130_fd_pr__cap_mim_m3_1_EN3Q86  sky130_fd_pr__cap_mim_m3_1_EN3Q86_0
timestamp 1662322327
transform 1 0 4943 0 1 3949
box -1750 -2240 1647 2240
use sky130_fd_pr__res_high_po_2p85_7J2RPB  sky130_fd_pr__res_high_po_2p85_7J2RPB_0
timestamp 1662230297
transform 0 1 4968 -1 0 1241
box -451 -1808 451 1808
<< labels >>
rlabel metal4 -820 5600 1820 5800 1 vdd
port 1 n
rlabel metal4 -5380 660 -3460 860 5 vss
port 2 s
rlabel metal1 -4685 710 -750 770 5 bias_0p7
rlabel metal2 3009 907 3356 1047 5 out
rlabel space -2958 2352 -2652 2432 3 in_p
rlabel space -3188 2172 -2652 2252 3 in_n
rlabel metal2 -2480 2590 -1740 2670 5 first_stage_out
rlabel space -4615 2259 -4025 2339 5 diffpair_source
rlabel metal3 -3832 2660 -3700 4300 7 ppair_gate
flabel metal2 -2752 2172 -2652 2252 0 FreeSans 1600 0 0 0 in_n
port 3 nsew
flabel metal2 -2752 2352 -2652 2432 0 FreeSans 1600 0 0 0 in_p
port 4 nsew
flabel metal2 301 2157 647 2289 0 FreeSans 1600 0 0 0 out
port 5 nsew
flabel metal1 -1324 594 -1276 766 0 FreeSans 1600 0 0 0 bias_0p7
port 6 nsew
<< end >>
