magic
tech sky130A
magscale 1 2
timestamp 1662519997
<< locali >>
rect 5840 10060 6580 10100
rect 7190 10060 7410 10100
rect 7990 10060 8210 10100
rect 8790 10060 9010 10100
rect 5840 9550 6590 9590
rect 7190 9540 7410 9580
rect 7990 9540 8210 9580
rect 8790 9540 9010 9580
<< metal1 >>
rect 5160 10000 5740 10040
rect 5160 9640 5200 10000
rect 5700 9640 5740 10000
rect 6570 10010 6640 10130
rect 7370 10010 7440 10130
rect 8170 10010 8240 10130
rect 8970 10010 9040 10130
rect 6570 9950 6980 10010
rect 7370 9950 7780 10010
rect 8170 9950 8580 10010
rect 8970 9950 9380 10010
rect 6570 9690 6640 9950
rect 6670 9910 6750 9920
rect 6670 9850 6680 9910
rect 6740 9850 6750 9910
rect 6670 9840 6750 9850
rect 6680 9720 6730 9840
rect 6780 9800 6830 9920
rect 6860 9910 6940 9920
rect 6860 9850 6870 9910
rect 6930 9850 6940 9910
rect 6860 9840 6940 9850
rect 6760 9790 6840 9800
rect 6760 9730 6770 9790
rect 6830 9730 6840 9790
rect 6760 9720 6840 9730
rect 6870 9720 6930 9840
rect 6970 9810 7030 9920
rect 7060 9910 7140 9920
rect 7060 9850 7070 9910
rect 7130 9850 7140 9910
rect 7060 9840 7140 9850
rect 7060 9830 7120 9840
rect 6960 9800 7030 9810
rect 6960 9790 7040 9800
rect 6960 9730 6970 9790
rect 7030 9730 7040 9790
rect 6960 9720 7040 9730
rect 7070 9720 7120 9830
rect 7370 9690 7440 9950
rect 7470 9910 7550 9920
rect 7470 9850 7480 9910
rect 7540 9850 7550 9910
rect 7470 9840 7550 9850
rect 7480 9720 7530 9840
rect 7580 9800 7630 9920
rect 7660 9910 7740 9920
rect 7660 9850 7670 9910
rect 7730 9850 7740 9910
rect 7660 9840 7740 9850
rect 7560 9790 7640 9800
rect 7560 9730 7570 9790
rect 7630 9730 7640 9790
rect 7560 9720 7640 9730
rect 7670 9720 7730 9840
rect 7770 9810 7830 9920
rect 7860 9910 7940 9920
rect 7860 9850 7870 9910
rect 7930 9850 7940 9910
rect 7860 9840 7940 9850
rect 7860 9830 7920 9840
rect 7760 9800 7830 9810
rect 7760 9790 7840 9800
rect 7760 9730 7770 9790
rect 7830 9730 7840 9790
rect 7760 9720 7840 9730
rect 7868 9720 7920 9830
rect 8170 9690 8240 9950
rect 8270 9910 8350 9920
rect 8270 9850 8280 9910
rect 8340 9850 8350 9910
rect 8270 9840 8350 9850
rect 8280 9720 8330 9840
rect 8380 9800 8430 9920
rect 8460 9910 8540 9920
rect 8460 9850 8470 9910
rect 8530 9850 8540 9910
rect 8460 9840 8540 9850
rect 8360 9790 8440 9800
rect 8360 9730 8370 9790
rect 8430 9730 8440 9790
rect 8360 9720 8440 9730
rect 8470 9720 8530 9840
rect 8570 9810 8630 9920
rect 8660 9910 8740 9920
rect 8660 9850 8670 9910
rect 8730 9850 8740 9910
rect 8660 9840 8740 9850
rect 8660 9830 8720 9840
rect 8560 9800 8630 9810
rect 8560 9790 8640 9800
rect 8560 9730 8570 9790
rect 8630 9730 8640 9790
rect 8560 9720 8640 9730
rect 8668 9720 8720 9830
rect 8970 9690 9040 9950
rect 9070 9910 9150 9920
rect 9070 9850 9080 9910
rect 9140 9850 9150 9910
rect 9070 9840 9150 9850
rect 9080 9720 9130 9840
rect 9180 9800 9230 9920
rect 9260 9910 9340 9920
rect 9260 9850 9270 9910
rect 9330 9850 9340 9910
rect 9260 9840 9340 9850
rect 9160 9790 9240 9800
rect 9160 9730 9170 9790
rect 9230 9730 9240 9790
rect 9160 9720 9240 9730
rect 9270 9720 9330 9840
rect 9370 9810 9430 9920
rect 9460 9910 9540 9920
rect 9460 9850 9470 9910
rect 9530 9850 9540 9910
rect 9460 9840 9540 9850
rect 9460 9830 9520 9840
rect 9360 9800 9430 9810
rect 9360 9790 9440 9800
rect 9360 9730 9370 9790
rect 9430 9730 9440 9790
rect 9360 9720 9440 9730
rect 9468 9720 9520 9830
rect 6570 9640 7080 9690
rect 7370 9640 7880 9690
rect 8170 9640 8680 9690
rect 8970 9640 9480 9690
rect 5160 9600 5740 9640
rect 5100 1200 5780 1240
rect 5100 740 5140 1200
rect 5740 740 5780 1200
rect 5100 700 5780 740
<< via1 >>
rect 5200 9640 5700 10000
rect 6680 9850 6740 9910
rect 6870 9850 6930 9910
rect 6770 9730 6830 9790
rect 7070 9850 7130 9910
rect 6970 9730 7030 9790
rect 7480 9850 7540 9910
rect 7670 9850 7730 9910
rect 7570 9730 7630 9790
rect 7870 9850 7930 9910
rect 7770 9730 7830 9790
rect 8280 9850 8340 9910
rect 8470 9850 8530 9910
rect 8370 9730 8430 9790
rect 8670 9850 8730 9910
rect 8570 9730 8630 9790
rect 9080 9850 9140 9910
rect 9270 9850 9330 9910
rect 9170 9730 9230 9790
rect 9470 9850 9530 9910
rect 9370 9730 9430 9790
rect 5140 740 5740 1200
<< metal2 >>
rect 7670 10040 7870 10060
rect 8470 10040 8670 10060
rect 9270 10040 9470 10060
rect 5160 10000 9540 10040
rect 5160 9640 5200 10000
rect 5700 9680 6080 10000
rect 6400 9910 9540 10000
rect 6400 9850 6680 9910
rect 6740 9850 6870 9910
rect 6930 9850 7070 9910
rect 7130 9850 7480 9910
rect 7540 9850 7670 9910
rect 7730 9850 7870 9910
rect 7930 9850 8280 9910
rect 8340 9850 8470 9910
rect 8530 9850 8670 9910
rect 8730 9850 9080 9910
rect 9140 9850 9270 9910
rect 9330 9850 9470 9910
rect 9530 9850 9540 9910
rect 6400 9840 9540 9850
rect 6400 9680 6440 9840
rect 5700 9640 6440 9680
rect 6540 9790 9570 9800
rect 6540 9730 6770 9790
rect 6830 9730 6970 9790
rect 7030 9730 7570 9790
rect 7630 9730 7770 9790
rect 7830 9730 8370 9790
rect 8430 9730 8570 9790
rect 8630 9730 9170 9790
rect 9230 9730 9370 9790
rect 9430 9730 9570 9790
rect 5160 9600 5740 9640
rect 6540 9510 9570 9730
rect 6540 9360 6830 9510
rect 5000 9070 6830 9360
rect 5000 1200 5780 1240
rect 5000 740 5140 1200
rect 5740 740 5780 1200
rect 5000 600 5780 740
<< via2 >>
rect 6080 9680 6400 10000
rect 5140 740 5740 1200
<< metal3 >>
rect 6040 10000 6440 10040
rect 6040 9680 6080 10000
rect 6400 9680 6440 10000
rect 6040 9640 6440 9680
rect 5100 1200 6040 1240
rect 5100 740 5140 1200
rect 5740 740 6040 1200
rect 5100 700 6040 740
<< via3 >>
rect 6080 9680 6400 10000
<< metal4 >>
rect 6040 10000 6440 10040
rect 6040 9680 6080 10000
rect 6400 9680 6440 10000
rect 6040 6420 6440 9680
rect 6040 590 6430 1670
use sky130_fd_pr__cap_mim_m3_1_4RCNTW  XC1
timestamp 1662404926
transform 1 0 8050 0 1 3700
box -2150 -3100 2149 3100
use sky130_fd_pr__nfet_01v8_lvt_HNLS5R  XM25 
timestamp 1662515274
transform 1 0 8499 0 -1 9820
box -359 -310 359 310
use sky130_fd_pr__nfet_01v8_lvt_HNLS5R  XM26
timestamp 1662515274
transform 1 0 9299 0 -1 9820
box -359 -310 359 310
use sky130_fd_pr__nfet_01v8_lvt_HNLS5R  XM27
timestamp 1662515274
transform 1 0 7699 0 -1 9820
box -359 -310 359 310
use sky130_fd_pr__nfet_01v8_lvt_HNLS5R  XM28
timestamp 1662515274
transform 1 0 6899 0 -1 9820
box -359 -310 359 310
use sky130_fd_pr__res_high_po_2p85_MXEQGY  XR18 
timestamp 1662404926
transform 1 0 5451 0 1 5398
box -451 -4798 451 4798
<< labels >>
rlabel metal2 5000 600 5140 1240 1 GND
rlabel metal1 6570 9950 6640 10130 1 IN1
rlabel metal2 5000 9070 6830 9360 1 VDD
rlabel metal1 7370 9640 7440 10130 1 IN2
rlabel metal1 8170 9640 8240 10130 1 IN3
rlabel metal1 8970 9640 9040 10130 1 IN4
rlabel metal4 6040 590 6430 1670 1 AMP
rlabel locali 5840 10060 6580 10100 1 SUB
<< end >>
