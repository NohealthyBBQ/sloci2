magic
tech sky130A
magscale 1 2
timestamp 1672264357
<< nwell >>
rect -2457 -3537 2457 3537
<< pmoslvt >>
rect -2261 118 -1861 3318
rect -1803 118 -1403 3318
rect -1345 118 -945 3318
rect -887 118 -487 3318
rect -429 118 -29 3318
rect 29 118 429 3318
rect 487 118 887 3318
rect 945 118 1345 3318
rect 1403 118 1803 3318
rect 1861 118 2261 3318
rect -2261 -3318 -1861 -118
rect -1803 -3318 -1403 -118
rect -1345 -3318 -945 -118
rect -887 -3318 -487 -118
rect -429 -3318 -29 -118
rect 29 -3318 429 -118
rect 487 -3318 887 -118
rect 945 -3318 1345 -118
rect 1403 -3318 1803 -118
rect 1861 -3318 2261 -118
<< pdiff >>
rect -2319 3306 -2261 3318
rect -2319 130 -2307 3306
rect -2273 130 -2261 3306
rect -2319 118 -2261 130
rect -1861 3306 -1803 3318
rect -1861 130 -1849 3306
rect -1815 130 -1803 3306
rect -1861 118 -1803 130
rect -1403 3306 -1345 3318
rect -1403 130 -1391 3306
rect -1357 130 -1345 3306
rect -1403 118 -1345 130
rect -945 3306 -887 3318
rect -945 130 -933 3306
rect -899 130 -887 3306
rect -945 118 -887 130
rect -487 3306 -429 3318
rect -487 130 -475 3306
rect -441 130 -429 3306
rect -487 118 -429 130
rect -29 3306 29 3318
rect -29 130 -17 3306
rect 17 130 29 3306
rect -29 118 29 130
rect 429 3306 487 3318
rect 429 130 441 3306
rect 475 130 487 3306
rect 429 118 487 130
rect 887 3306 945 3318
rect 887 130 899 3306
rect 933 130 945 3306
rect 887 118 945 130
rect 1345 3306 1403 3318
rect 1345 130 1357 3306
rect 1391 130 1403 3306
rect 1345 118 1403 130
rect 1803 3306 1861 3318
rect 1803 130 1815 3306
rect 1849 130 1861 3306
rect 1803 118 1861 130
rect 2261 3306 2319 3318
rect 2261 130 2273 3306
rect 2307 130 2319 3306
rect 2261 118 2319 130
rect -2319 -130 -2261 -118
rect -2319 -3306 -2307 -130
rect -2273 -3306 -2261 -130
rect -2319 -3318 -2261 -3306
rect -1861 -130 -1803 -118
rect -1861 -3306 -1849 -130
rect -1815 -3306 -1803 -130
rect -1861 -3318 -1803 -3306
rect -1403 -130 -1345 -118
rect -1403 -3306 -1391 -130
rect -1357 -3306 -1345 -130
rect -1403 -3318 -1345 -3306
rect -945 -130 -887 -118
rect -945 -3306 -933 -130
rect -899 -3306 -887 -130
rect -945 -3318 -887 -3306
rect -487 -130 -429 -118
rect -487 -3306 -475 -130
rect -441 -3306 -429 -130
rect -487 -3318 -429 -3306
rect -29 -130 29 -118
rect -29 -3306 -17 -130
rect 17 -3306 29 -130
rect -29 -3318 29 -3306
rect 429 -130 487 -118
rect 429 -3306 441 -130
rect 475 -3306 487 -130
rect 429 -3318 487 -3306
rect 887 -130 945 -118
rect 887 -3306 899 -130
rect 933 -3306 945 -130
rect 887 -3318 945 -3306
rect 1345 -130 1403 -118
rect 1345 -3306 1357 -130
rect 1391 -3306 1403 -130
rect 1345 -3318 1403 -3306
rect 1803 -130 1861 -118
rect 1803 -3306 1815 -130
rect 1849 -3306 1861 -130
rect 1803 -3318 1861 -3306
rect 2261 -130 2319 -118
rect 2261 -3306 2273 -130
rect 2307 -3306 2319 -130
rect 2261 -3318 2319 -3306
<< pdiffc >>
rect -2307 130 -2273 3306
rect -1849 130 -1815 3306
rect -1391 130 -1357 3306
rect -933 130 -899 3306
rect -475 130 -441 3306
rect -17 130 17 3306
rect 441 130 475 3306
rect 899 130 933 3306
rect 1357 130 1391 3306
rect 1815 130 1849 3306
rect 2273 130 2307 3306
rect -2307 -3306 -2273 -130
rect -1849 -3306 -1815 -130
rect -1391 -3306 -1357 -130
rect -933 -3306 -899 -130
rect -475 -3306 -441 -130
rect -17 -3306 17 -130
rect 441 -3306 475 -130
rect 899 -3306 933 -130
rect 1357 -3306 1391 -130
rect 1815 -3306 1849 -130
rect 2273 -3306 2307 -130
<< nsubdiff >>
rect -2421 3467 -2325 3501
rect 2325 3467 2421 3501
rect -2421 3405 -2387 3467
rect 2387 3405 2421 3467
rect -2421 -3467 -2387 -3405
rect 2387 -3467 2421 -3405
rect -2421 -3501 -2325 -3467
rect 2325 -3501 2421 -3467
<< nsubdiffcont >>
rect -2325 3467 2325 3501
rect -2421 -3405 -2387 3405
rect 2387 -3405 2421 3405
rect -2325 -3501 2325 -3467
<< poly >>
rect -2261 3399 -1861 3415
rect -2261 3365 -2245 3399
rect -1877 3365 -1861 3399
rect -2261 3318 -1861 3365
rect -1803 3399 -1403 3415
rect -1803 3365 -1787 3399
rect -1419 3365 -1403 3399
rect -1803 3318 -1403 3365
rect -1345 3399 -945 3415
rect -1345 3365 -1329 3399
rect -961 3365 -945 3399
rect -1345 3318 -945 3365
rect -887 3399 -487 3415
rect -887 3365 -871 3399
rect -503 3365 -487 3399
rect -887 3318 -487 3365
rect -429 3399 -29 3415
rect -429 3365 -413 3399
rect -45 3365 -29 3399
rect -429 3318 -29 3365
rect 29 3399 429 3415
rect 29 3365 45 3399
rect 413 3365 429 3399
rect 29 3318 429 3365
rect 487 3399 887 3415
rect 487 3365 503 3399
rect 871 3365 887 3399
rect 487 3318 887 3365
rect 945 3399 1345 3415
rect 945 3365 961 3399
rect 1329 3365 1345 3399
rect 945 3318 1345 3365
rect 1403 3399 1803 3415
rect 1403 3365 1419 3399
rect 1787 3365 1803 3399
rect 1403 3318 1803 3365
rect 1861 3399 2261 3415
rect 1861 3365 1877 3399
rect 2245 3365 2261 3399
rect 1861 3318 2261 3365
rect -2261 71 -1861 118
rect -2261 37 -2245 71
rect -1877 37 -1861 71
rect -2261 21 -1861 37
rect -1803 71 -1403 118
rect -1803 37 -1787 71
rect -1419 37 -1403 71
rect -1803 21 -1403 37
rect -1345 71 -945 118
rect -1345 37 -1329 71
rect -961 37 -945 71
rect -1345 21 -945 37
rect -887 71 -487 118
rect -887 37 -871 71
rect -503 37 -487 71
rect -887 21 -487 37
rect -429 71 -29 118
rect -429 37 -413 71
rect -45 37 -29 71
rect -429 21 -29 37
rect 29 71 429 118
rect 29 37 45 71
rect 413 37 429 71
rect 29 21 429 37
rect 487 71 887 118
rect 487 37 503 71
rect 871 37 887 71
rect 487 21 887 37
rect 945 71 1345 118
rect 945 37 961 71
rect 1329 37 1345 71
rect 945 21 1345 37
rect 1403 71 1803 118
rect 1403 37 1419 71
rect 1787 37 1803 71
rect 1403 21 1803 37
rect 1861 71 2261 118
rect 1861 37 1877 71
rect 2245 37 2261 71
rect 1861 21 2261 37
rect -2261 -37 -1861 -21
rect -2261 -71 -2245 -37
rect -1877 -71 -1861 -37
rect -2261 -118 -1861 -71
rect -1803 -37 -1403 -21
rect -1803 -71 -1787 -37
rect -1419 -71 -1403 -37
rect -1803 -118 -1403 -71
rect -1345 -37 -945 -21
rect -1345 -71 -1329 -37
rect -961 -71 -945 -37
rect -1345 -118 -945 -71
rect -887 -37 -487 -21
rect -887 -71 -871 -37
rect -503 -71 -487 -37
rect -887 -118 -487 -71
rect -429 -37 -29 -21
rect -429 -71 -413 -37
rect -45 -71 -29 -37
rect -429 -118 -29 -71
rect 29 -37 429 -21
rect 29 -71 45 -37
rect 413 -71 429 -37
rect 29 -118 429 -71
rect 487 -37 887 -21
rect 487 -71 503 -37
rect 871 -71 887 -37
rect 487 -118 887 -71
rect 945 -37 1345 -21
rect 945 -71 961 -37
rect 1329 -71 1345 -37
rect 945 -118 1345 -71
rect 1403 -37 1803 -21
rect 1403 -71 1419 -37
rect 1787 -71 1803 -37
rect 1403 -118 1803 -71
rect 1861 -37 2261 -21
rect 1861 -71 1877 -37
rect 2245 -71 2261 -37
rect 1861 -118 2261 -71
rect -2261 -3365 -1861 -3318
rect -2261 -3399 -2245 -3365
rect -1877 -3399 -1861 -3365
rect -2261 -3415 -1861 -3399
rect -1803 -3365 -1403 -3318
rect -1803 -3399 -1787 -3365
rect -1419 -3399 -1403 -3365
rect -1803 -3415 -1403 -3399
rect -1345 -3365 -945 -3318
rect -1345 -3399 -1329 -3365
rect -961 -3399 -945 -3365
rect -1345 -3415 -945 -3399
rect -887 -3365 -487 -3318
rect -887 -3399 -871 -3365
rect -503 -3399 -487 -3365
rect -887 -3415 -487 -3399
rect -429 -3365 -29 -3318
rect -429 -3399 -413 -3365
rect -45 -3399 -29 -3365
rect -429 -3415 -29 -3399
rect 29 -3365 429 -3318
rect 29 -3399 45 -3365
rect 413 -3399 429 -3365
rect 29 -3415 429 -3399
rect 487 -3365 887 -3318
rect 487 -3399 503 -3365
rect 871 -3399 887 -3365
rect 487 -3415 887 -3399
rect 945 -3365 1345 -3318
rect 945 -3399 961 -3365
rect 1329 -3399 1345 -3365
rect 945 -3415 1345 -3399
rect 1403 -3365 1803 -3318
rect 1403 -3399 1419 -3365
rect 1787 -3399 1803 -3365
rect 1403 -3415 1803 -3399
rect 1861 -3365 2261 -3318
rect 1861 -3399 1877 -3365
rect 2245 -3399 2261 -3365
rect 1861 -3415 2261 -3399
<< polycont >>
rect -2245 3365 -1877 3399
rect -1787 3365 -1419 3399
rect -1329 3365 -961 3399
rect -871 3365 -503 3399
rect -413 3365 -45 3399
rect 45 3365 413 3399
rect 503 3365 871 3399
rect 961 3365 1329 3399
rect 1419 3365 1787 3399
rect 1877 3365 2245 3399
rect -2245 37 -1877 71
rect -1787 37 -1419 71
rect -1329 37 -961 71
rect -871 37 -503 71
rect -413 37 -45 71
rect 45 37 413 71
rect 503 37 871 71
rect 961 37 1329 71
rect 1419 37 1787 71
rect 1877 37 2245 71
rect -2245 -71 -1877 -37
rect -1787 -71 -1419 -37
rect -1329 -71 -961 -37
rect -871 -71 -503 -37
rect -413 -71 -45 -37
rect 45 -71 413 -37
rect 503 -71 871 -37
rect 961 -71 1329 -37
rect 1419 -71 1787 -37
rect 1877 -71 2245 -37
rect -2245 -3399 -1877 -3365
rect -1787 -3399 -1419 -3365
rect -1329 -3399 -961 -3365
rect -871 -3399 -503 -3365
rect -413 -3399 -45 -3365
rect 45 -3399 413 -3365
rect 503 -3399 871 -3365
rect 961 -3399 1329 -3365
rect 1419 -3399 1787 -3365
rect 1877 -3399 2245 -3365
<< locali >>
rect -2421 3467 -2325 3501
rect 2325 3467 2421 3501
rect -2421 3405 -2387 3467
rect 2387 3405 2421 3467
rect -2261 3365 -2245 3399
rect -1877 3365 -1861 3399
rect -1803 3365 -1787 3399
rect -1419 3365 -1403 3399
rect -1345 3365 -1329 3399
rect -961 3365 -945 3399
rect -887 3365 -871 3399
rect -503 3365 -487 3399
rect -429 3365 -413 3399
rect -45 3365 -29 3399
rect 29 3365 45 3399
rect 413 3365 429 3399
rect 487 3365 503 3399
rect 871 3365 887 3399
rect 945 3365 961 3399
rect 1329 3365 1345 3399
rect 1403 3365 1419 3399
rect 1787 3365 1803 3399
rect 1861 3365 1877 3399
rect 2245 3365 2261 3399
rect -2307 3306 -2273 3322
rect -2307 114 -2273 130
rect -1849 3306 -1815 3322
rect -1849 114 -1815 130
rect -1391 3306 -1357 3322
rect -1391 114 -1357 130
rect -933 3306 -899 3322
rect -933 114 -899 130
rect -475 3306 -441 3322
rect -475 114 -441 130
rect -17 3306 17 3322
rect -17 114 17 130
rect 441 3306 475 3322
rect 441 114 475 130
rect 899 3306 933 3322
rect 899 114 933 130
rect 1357 3306 1391 3322
rect 1357 114 1391 130
rect 1815 3306 1849 3322
rect 1815 114 1849 130
rect 2273 3306 2307 3322
rect 2273 114 2307 130
rect -2261 37 -2245 71
rect -1877 37 -1861 71
rect -1803 37 -1787 71
rect -1419 37 -1403 71
rect -1345 37 -1329 71
rect -961 37 -945 71
rect -887 37 -871 71
rect -503 37 -487 71
rect -429 37 -413 71
rect -45 37 -29 71
rect 29 37 45 71
rect 413 37 429 71
rect 487 37 503 71
rect 871 37 887 71
rect 945 37 961 71
rect 1329 37 1345 71
rect 1403 37 1419 71
rect 1787 37 1803 71
rect 1861 37 1877 71
rect 2245 37 2261 71
rect -2261 -71 -2245 -37
rect -1877 -71 -1861 -37
rect -1803 -71 -1787 -37
rect -1419 -71 -1403 -37
rect -1345 -71 -1329 -37
rect -961 -71 -945 -37
rect -887 -71 -871 -37
rect -503 -71 -487 -37
rect -429 -71 -413 -37
rect -45 -71 -29 -37
rect 29 -71 45 -37
rect 413 -71 429 -37
rect 487 -71 503 -37
rect 871 -71 887 -37
rect 945 -71 961 -37
rect 1329 -71 1345 -37
rect 1403 -71 1419 -37
rect 1787 -71 1803 -37
rect 1861 -71 1877 -37
rect 2245 -71 2261 -37
rect -2307 -130 -2273 -114
rect -2307 -3322 -2273 -3306
rect -1849 -130 -1815 -114
rect -1849 -3322 -1815 -3306
rect -1391 -130 -1357 -114
rect -1391 -3322 -1357 -3306
rect -933 -130 -899 -114
rect -933 -3322 -899 -3306
rect -475 -130 -441 -114
rect -475 -3322 -441 -3306
rect -17 -130 17 -114
rect -17 -3322 17 -3306
rect 441 -130 475 -114
rect 441 -3322 475 -3306
rect 899 -130 933 -114
rect 899 -3322 933 -3306
rect 1357 -130 1391 -114
rect 1357 -3322 1391 -3306
rect 1815 -130 1849 -114
rect 1815 -3322 1849 -3306
rect 2273 -130 2307 -114
rect 2273 -3322 2307 -3306
rect -2261 -3399 -2245 -3365
rect -1877 -3399 -1861 -3365
rect -1803 -3399 -1787 -3365
rect -1419 -3399 -1403 -3365
rect -1345 -3399 -1329 -3365
rect -961 -3399 -945 -3365
rect -887 -3399 -871 -3365
rect -503 -3399 -487 -3365
rect -429 -3399 -413 -3365
rect -45 -3399 -29 -3365
rect 29 -3399 45 -3365
rect 413 -3399 429 -3365
rect 487 -3399 503 -3365
rect 871 -3399 887 -3365
rect 945 -3399 961 -3365
rect 1329 -3399 1345 -3365
rect 1403 -3399 1419 -3365
rect 1787 -3399 1803 -3365
rect 1861 -3399 1877 -3365
rect 2245 -3399 2261 -3365
rect -2421 -3467 -2387 -3405
rect 2387 -3467 2421 -3405
rect -2421 -3501 -2325 -3467
rect 2325 -3501 2421 -3467
<< viali >>
rect -2245 3365 -1877 3399
rect -1787 3365 -1419 3399
rect -1329 3365 -961 3399
rect -871 3365 -503 3399
rect -413 3365 -45 3399
rect 45 3365 413 3399
rect 503 3365 871 3399
rect 961 3365 1329 3399
rect 1419 3365 1787 3399
rect 1877 3365 2245 3399
rect -2307 130 -2273 3306
rect -1849 130 -1815 3306
rect -1391 130 -1357 3306
rect -933 130 -899 3306
rect -475 130 -441 3306
rect -17 130 17 3306
rect 441 130 475 3306
rect 899 130 933 3306
rect 1357 130 1391 3306
rect 1815 130 1849 3306
rect 2273 130 2307 3306
rect -2245 37 -1877 71
rect -1787 37 -1419 71
rect -1329 37 -961 71
rect -871 37 -503 71
rect -413 37 -45 71
rect 45 37 413 71
rect 503 37 871 71
rect 961 37 1329 71
rect 1419 37 1787 71
rect 1877 37 2245 71
rect -2245 -71 -1877 -37
rect -1787 -71 -1419 -37
rect -1329 -71 -961 -37
rect -871 -71 -503 -37
rect -413 -71 -45 -37
rect 45 -71 413 -37
rect 503 -71 871 -37
rect 961 -71 1329 -37
rect 1419 -71 1787 -37
rect 1877 -71 2245 -37
rect -2307 -3306 -2273 -130
rect -1849 -3306 -1815 -130
rect -1391 -3306 -1357 -130
rect -933 -3306 -899 -130
rect -475 -3306 -441 -130
rect -17 -3306 17 -130
rect 441 -3306 475 -130
rect 899 -3306 933 -130
rect 1357 -3306 1391 -130
rect 1815 -3306 1849 -130
rect 2273 -3306 2307 -130
rect -2245 -3399 -1877 -3365
rect -1787 -3399 -1419 -3365
rect -1329 -3399 -961 -3365
rect -871 -3399 -503 -3365
rect -413 -3399 -45 -3365
rect 45 -3399 413 -3365
rect 503 -3399 871 -3365
rect 961 -3399 1329 -3365
rect 1419 -3399 1787 -3365
rect 1877 -3399 2245 -3365
<< metal1 >>
rect -2257 3399 -1865 3405
rect -2257 3365 -2245 3399
rect -1877 3365 -1865 3399
rect -2257 3359 -1865 3365
rect -1799 3399 -1407 3405
rect -1799 3365 -1787 3399
rect -1419 3365 -1407 3399
rect -1799 3359 -1407 3365
rect -1341 3399 -949 3405
rect -1341 3365 -1329 3399
rect -961 3365 -949 3399
rect -1341 3359 -949 3365
rect -883 3399 -491 3405
rect -883 3365 -871 3399
rect -503 3365 -491 3399
rect -883 3359 -491 3365
rect -425 3399 -33 3405
rect -425 3365 -413 3399
rect -45 3365 -33 3399
rect -425 3359 -33 3365
rect 33 3399 425 3405
rect 33 3365 45 3399
rect 413 3365 425 3399
rect 33 3359 425 3365
rect 491 3399 883 3405
rect 491 3365 503 3399
rect 871 3365 883 3399
rect 491 3359 883 3365
rect 949 3399 1341 3405
rect 949 3365 961 3399
rect 1329 3365 1341 3399
rect 949 3359 1341 3365
rect 1407 3399 1799 3405
rect 1407 3365 1419 3399
rect 1787 3365 1799 3399
rect 1407 3359 1799 3365
rect 1865 3399 2257 3405
rect 1865 3365 1877 3399
rect 2245 3365 2257 3399
rect 1865 3359 2257 3365
rect -2313 3306 -2267 3318
rect -2313 130 -2307 3306
rect -2273 130 -2267 3306
rect -2313 118 -2267 130
rect -1855 3306 -1809 3318
rect -1855 130 -1849 3306
rect -1815 130 -1809 3306
rect -1855 118 -1809 130
rect -1397 3306 -1351 3318
rect -1397 130 -1391 3306
rect -1357 130 -1351 3306
rect -1397 118 -1351 130
rect -939 3306 -893 3318
rect -939 130 -933 3306
rect -899 130 -893 3306
rect -939 118 -893 130
rect -481 3306 -435 3318
rect -481 130 -475 3306
rect -441 130 -435 3306
rect -481 118 -435 130
rect -23 3306 23 3318
rect -23 130 -17 3306
rect 17 130 23 3306
rect -23 118 23 130
rect 435 3306 481 3318
rect 435 130 441 3306
rect 475 130 481 3306
rect 435 118 481 130
rect 893 3306 939 3318
rect 893 130 899 3306
rect 933 130 939 3306
rect 893 118 939 130
rect 1351 3306 1397 3318
rect 1351 130 1357 3306
rect 1391 130 1397 3306
rect 1351 118 1397 130
rect 1809 3306 1855 3318
rect 1809 130 1815 3306
rect 1849 130 1855 3306
rect 1809 118 1855 130
rect 2267 3306 2313 3318
rect 2267 130 2273 3306
rect 2307 130 2313 3306
rect 2267 118 2313 130
rect -2257 71 -1865 77
rect -2257 37 -2245 71
rect -1877 37 -1865 71
rect -2257 31 -1865 37
rect -1799 71 -1407 77
rect -1799 37 -1787 71
rect -1419 37 -1407 71
rect -1799 31 -1407 37
rect -1341 71 -949 77
rect -1341 37 -1329 71
rect -961 37 -949 71
rect -1341 31 -949 37
rect -883 71 -491 77
rect -883 37 -871 71
rect -503 37 -491 71
rect -883 31 -491 37
rect -425 71 -33 77
rect -425 37 -413 71
rect -45 37 -33 71
rect -425 31 -33 37
rect 33 71 425 77
rect 33 37 45 71
rect 413 37 425 71
rect 33 31 425 37
rect 491 71 883 77
rect 491 37 503 71
rect 871 37 883 71
rect 491 31 883 37
rect 949 71 1341 77
rect 949 37 961 71
rect 1329 37 1341 71
rect 949 31 1341 37
rect 1407 71 1799 77
rect 1407 37 1419 71
rect 1787 37 1799 71
rect 1407 31 1799 37
rect 1865 71 2257 77
rect 1865 37 1877 71
rect 2245 37 2257 71
rect 1865 31 2257 37
rect -2257 -37 -1865 -31
rect -2257 -71 -2245 -37
rect -1877 -71 -1865 -37
rect -2257 -77 -1865 -71
rect -1799 -37 -1407 -31
rect -1799 -71 -1787 -37
rect -1419 -71 -1407 -37
rect -1799 -77 -1407 -71
rect -1341 -37 -949 -31
rect -1341 -71 -1329 -37
rect -961 -71 -949 -37
rect -1341 -77 -949 -71
rect -883 -37 -491 -31
rect -883 -71 -871 -37
rect -503 -71 -491 -37
rect -883 -77 -491 -71
rect -425 -37 -33 -31
rect -425 -71 -413 -37
rect -45 -71 -33 -37
rect -425 -77 -33 -71
rect 33 -37 425 -31
rect 33 -71 45 -37
rect 413 -71 425 -37
rect 33 -77 425 -71
rect 491 -37 883 -31
rect 491 -71 503 -37
rect 871 -71 883 -37
rect 491 -77 883 -71
rect 949 -37 1341 -31
rect 949 -71 961 -37
rect 1329 -71 1341 -37
rect 949 -77 1341 -71
rect 1407 -37 1799 -31
rect 1407 -71 1419 -37
rect 1787 -71 1799 -37
rect 1407 -77 1799 -71
rect 1865 -37 2257 -31
rect 1865 -71 1877 -37
rect 2245 -71 2257 -37
rect 1865 -77 2257 -71
rect -2313 -130 -2267 -118
rect -2313 -3306 -2307 -130
rect -2273 -3306 -2267 -130
rect -2313 -3318 -2267 -3306
rect -1855 -130 -1809 -118
rect -1855 -3306 -1849 -130
rect -1815 -3306 -1809 -130
rect -1855 -3318 -1809 -3306
rect -1397 -130 -1351 -118
rect -1397 -3306 -1391 -130
rect -1357 -3306 -1351 -130
rect -1397 -3318 -1351 -3306
rect -939 -130 -893 -118
rect -939 -3306 -933 -130
rect -899 -3306 -893 -130
rect -939 -3318 -893 -3306
rect -481 -130 -435 -118
rect -481 -3306 -475 -130
rect -441 -3306 -435 -130
rect -481 -3318 -435 -3306
rect -23 -130 23 -118
rect -23 -3306 -17 -130
rect 17 -3306 23 -130
rect -23 -3318 23 -3306
rect 435 -130 481 -118
rect 435 -3306 441 -130
rect 475 -3306 481 -130
rect 435 -3318 481 -3306
rect 893 -130 939 -118
rect 893 -3306 899 -130
rect 933 -3306 939 -130
rect 893 -3318 939 -3306
rect 1351 -130 1397 -118
rect 1351 -3306 1357 -130
rect 1391 -3306 1397 -130
rect 1351 -3318 1397 -3306
rect 1809 -130 1855 -118
rect 1809 -3306 1815 -130
rect 1849 -3306 1855 -130
rect 1809 -3318 1855 -3306
rect 2267 -130 2313 -118
rect 2267 -3306 2273 -130
rect 2307 -3306 2313 -130
rect 2267 -3318 2313 -3306
rect -2257 -3365 -1865 -3359
rect -2257 -3399 -2245 -3365
rect -1877 -3399 -1865 -3365
rect -2257 -3405 -1865 -3399
rect -1799 -3365 -1407 -3359
rect -1799 -3399 -1787 -3365
rect -1419 -3399 -1407 -3365
rect -1799 -3405 -1407 -3399
rect -1341 -3365 -949 -3359
rect -1341 -3399 -1329 -3365
rect -961 -3399 -949 -3365
rect -1341 -3405 -949 -3399
rect -883 -3365 -491 -3359
rect -883 -3399 -871 -3365
rect -503 -3399 -491 -3365
rect -883 -3405 -491 -3399
rect -425 -3365 -33 -3359
rect -425 -3399 -413 -3365
rect -45 -3399 -33 -3365
rect -425 -3405 -33 -3399
rect 33 -3365 425 -3359
rect 33 -3399 45 -3365
rect 413 -3399 425 -3365
rect 33 -3405 425 -3399
rect 491 -3365 883 -3359
rect 491 -3399 503 -3365
rect 871 -3399 883 -3365
rect 491 -3405 883 -3399
rect 949 -3365 1341 -3359
rect 949 -3399 961 -3365
rect 1329 -3399 1341 -3365
rect 949 -3405 1341 -3399
rect 1407 -3365 1799 -3359
rect 1407 -3399 1419 -3365
rect 1787 -3399 1799 -3365
rect 1407 -3405 1799 -3399
rect 1865 -3365 2257 -3359
rect 1865 -3399 1877 -3365
rect 2245 -3399 2257 -3365
rect 1865 -3405 2257 -3399
<< properties >>
string FIXED_BBOX -2404 -3484 2404 3484
string gencell sky130_fd_pr__pfet_01v8_lvt
string library sky130
string parameters w 16 l 2 m 2 nf 10 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.35 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
