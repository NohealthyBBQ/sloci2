magic
tech sky130A
magscale 1 2
timestamp 1672531254
<< metal4 >>
rect -200 50 200 107
rect -200 -107 200 -50
<< rmetal4 >>
rect -200 -50 200 50
<< properties >>
string gencell sky130_fd_pr__res_generic_m4
string library sky130
string parameters w 2 l 0.5 m 1 nx 1 wmin 0.30 lmin 0.30 rho 0.047 val 11.75m dummy 0 dw 0.0 term 0.0 roverlap 0
<< end >>
