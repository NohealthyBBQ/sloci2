magic
tech sky130A
timestamp 1672090903
<< pwell >>
rect -300 -155 299 155
<< nmoslvt >>
rect -200 -50 -185 50
rect -152 -50 -137 50
rect -104 -50 -89 50
rect -56 -50 -41 50
rect -8 -50 7 50
rect 40 -50 55 50
rect 88 -50 103 50
rect 136 -50 151 50
rect 184 -50 199 50
<< ndiff >>
rect -231 44 -200 50
rect -231 -44 -225 44
rect -208 -44 -200 44
rect -231 -50 -200 -44
rect -185 44 -152 50
rect -185 -44 -177 44
rect -160 -44 -152 44
rect -185 -50 -152 -44
rect -137 44 -104 50
rect -137 -44 -129 44
rect -112 -44 -104 44
rect -137 -50 -104 -44
rect -89 44 -56 50
rect -89 -44 -81 44
rect -64 -44 -56 44
rect -89 -50 -56 -44
rect -41 44 -8 50
rect -41 -44 -33 44
rect -16 -44 -8 44
rect -41 -50 -8 -44
rect 7 44 40 50
rect 7 -44 15 44
rect 32 -44 40 44
rect 7 -50 40 -44
rect 55 44 88 50
rect 55 -44 63 44
rect 80 -44 88 44
rect 55 -50 88 -44
rect 103 44 136 50
rect 103 -44 111 44
rect 128 -44 136 44
rect 103 -50 136 -44
rect 151 44 184 50
rect 151 -44 159 44
rect 176 -44 184 44
rect 151 -50 184 -44
rect 199 44 230 50
rect 199 -44 207 44
rect 224 -44 230 44
rect 199 -50 230 -44
<< ndiffc >>
rect -225 -44 -208 44
rect -177 -44 -160 44
rect -129 -44 -112 44
rect -81 -44 -64 44
rect -33 -44 -16 44
rect 15 -44 32 44
rect 63 -44 80 44
rect 111 -44 128 44
rect 159 -44 176 44
rect 207 -44 224 44
<< psubdiff >>
rect -282 120 -234 137
rect 233 120 281 137
rect -282 89 -265 120
rect 264 89 281 120
rect -282 -120 -265 -89
rect 264 -120 281 -89
rect -282 -137 -234 -120
rect 233 -137 281 -120
<< psubdiffcont >>
rect -234 120 233 137
rect -282 -89 -265 89
rect 264 -89 281 89
rect -234 -137 233 -120
<< poly >>
rect -200 50 -185 63
rect -152 50 -137 63
rect -104 50 -89 63
rect -56 50 -41 63
rect -8 50 7 63
rect 40 50 55 63
rect 88 50 103 63
rect 136 50 151 63
rect 184 50 199 63
rect -200 -61 -185 -50
rect -152 -61 -137 -50
rect -104 -61 -89 -50
rect -56 -61 -41 -50
rect -8 -61 7 -50
rect 40 -61 55 -50
rect 88 -61 103 -50
rect 136 -61 151 -50
rect 184 -61 199 -50
rect -209 -69 208 -61
rect -209 -86 183 -69
rect 200 -86 208 -69
rect 175 -94 208 -86
<< polycont >>
rect 183 -86 200 -69
<< locali >>
rect -282 120 -234 137
rect 233 120 281 137
rect -282 89 -265 120
rect 264 89 281 120
rect -225 44 -208 52
rect -225 -52 -208 -44
rect -177 44 -160 52
rect -177 -52 -160 -44
rect -129 44 -112 52
rect -129 -52 -112 -44
rect -81 44 -64 52
rect -81 -52 -64 -44
rect -33 44 -16 52
rect -33 -52 -16 -44
rect 15 44 32 52
rect 15 -52 32 -44
rect 63 44 80 52
rect 63 -52 80 -44
rect 111 44 128 52
rect 111 -52 128 -44
rect 159 44 176 52
rect 159 -52 176 -44
rect 207 44 224 52
rect 207 -52 224 -44
rect 175 -86 183 -69
rect 200 -86 208 -69
rect -282 -120 -265 -89
rect 264 -120 281 -89
rect -282 -137 -234 -120
rect 233 -137 281 -120
<< viali >>
rect -225 -44 -208 44
rect -177 -44 -160 44
rect -129 -44 -112 44
rect -81 -44 -64 44
rect -33 -44 -16 44
rect 15 -44 32 44
rect 63 -44 80 44
rect 111 -44 128 44
rect 159 -44 176 44
rect 207 -44 224 44
rect 183 -86 200 -69
<< metal1 >>
rect -228 44 -205 50
rect -228 -14 -225 44
rect -233 -17 -225 -14
rect -208 -14 -205 44
rect -185 47 -152 50
rect -185 17 -182 47
rect -155 17 -152 47
rect -185 14 -177 17
rect -208 -17 -200 -14
rect -233 -47 -230 -17
rect -203 -47 -200 -17
rect -233 -50 -200 -47
rect -180 -44 -177 14
rect -160 14 -152 17
rect -132 44 -109 50
rect -160 -44 -157 14
rect -132 -14 -129 44
rect -180 -50 -157 -44
rect -137 -17 -129 -14
rect -112 -14 -109 44
rect -89 47 -56 50
rect -89 17 -86 47
rect -59 17 -56 47
rect -89 14 -81 17
rect -112 -17 -104 -14
rect -137 -47 -134 -17
rect -107 -47 -104 -17
rect -137 -50 -104 -47
rect -84 -44 -81 14
rect -64 14 -56 17
rect -36 44 -13 50
rect -64 -44 -61 14
rect -36 -14 -33 44
rect -84 -50 -61 -44
rect -41 -17 -33 -14
rect -16 -14 -13 44
rect 7 47 40 50
rect 7 17 10 47
rect 37 17 40 47
rect 7 14 15 17
rect -16 -17 -8 -14
rect -41 -47 -38 -17
rect -11 -47 -8 -17
rect -41 -50 -8 -47
rect 12 -44 15 14
rect 32 14 40 17
rect 60 44 83 50
rect 32 -44 35 14
rect 60 -14 63 44
rect 12 -50 35 -44
rect 55 -17 63 -14
rect 80 -14 83 44
rect 103 47 136 50
rect 103 17 106 47
rect 133 17 136 47
rect 103 14 111 17
rect 80 -17 88 -14
rect 55 -47 58 -17
rect 85 -47 88 -17
rect 55 -50 88 -47
rect 108 -44 111 14
rect 128 14 136 17
rect 156 44 179 50
rect 128 -44 131 14
rect 156 -14 159 44
rect 108 -50 131 -44
rect 151 -17 159 -14
rect 176 -14 179 44
rect 199 47 232 50
rect 199 17 202 47
rect 229 17 232 47
rect 199 14 207 17
rect 176 -17 184 -14
rect 151 -47 154 -17
rect 181 -47 184 -17
rect 151 -50 184 -47
rect 204 -44 207 14
rect 224 14 232 17
rect 224 -44 227 14
rect 204 -50 227 -44
rect 175 -69 216 -66
rect 175 -86 183 -69
rect 200 -86 216 -69
rect 175 -94 216 -86
<< via1 >>
rect -182 44 -155 47
rect -182 17 -177 44
rect -177 17 -160 44
rect -160 17 -155 44
rect -230 -44 -225 -17
rect -225 -44 -208 -17
rect -208 -44 -203 -17
rect -230 -47 -203 -44
rect -86 44 -59 47
rect -86 17 -81 44
rect -81 17 -64 44
rect -64 17 -59 44
rect -134 -44 -129 -17
rect -129 -44 -112 -17
rect -112 -44 -107 -17
rect -134 -47 -107 -44
rect 10 44 37 47
rect 10 17 15 44
rect 15 17 32 44
rect 32 17 37 44
rect -38 -44 -33 -17
rect -33 -44 -16 -17
rect -16 -44 -11 -17
rect -38 -47 -11 -44
rect 106 44 133 47
rect 106 17 111 44
rect 111 17 128 44
rect 128 17 133 44
rect 58 -44 63 -17
rect 63 -44 80 -17
rect 80 -44 85 -17
rect 58 -47 85 -44
rect 202 44 229 47
rect 202 17 207 44
rect 207 17 224 44
rect 224 17 229 44
rect 154 -44 159 -17
rect 159 -44 176 -17
rect 176 -44 181 -17
rect 154 -47 181 -44
<< metal2 >>
rect -233 47 232 50
rect -233 17 -182 47
rect -155 17 -86 47
rect -59 17 10 47
rect 37 17 106 47
rect 133 17 202 47
rect 229 17 232 47
rect -233 14 232 17
rect -233 -17 230 -14
rect -233 -47 -230 -17
rect -203 -47 -134 -17
rect -107 -47 -38 -17
rect -11 -47 58 -17
rect 85 -47 154 -17
rect 181 -47 230 -17
rect -233 -50 230 -47
<< properties >>
string FIXED_BBOX -273 -128 273 128
string gencell sky130_fd_pr__nfet_01v8_lvt
string library sky130
string parameters w 1.0 l 0.15 m 1 nf 9 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
