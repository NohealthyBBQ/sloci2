magic
tech sky130A
magscale 1 2
timestamp 1662302892
<< pwell >>
rect -625 -1491 625 1491
<< nmoslvt >>
rect -429 943 -29 1343
rect 29 943 429 1343
rect -429 387 -29 787
rect 29 387 429 787
rect -429 -169 -29 231
rect 29 -169 429 231
rect -429 -725 -29 -325
rect 29 -725 429 -325
rect -429 -1281 -29 -881
rect 29 -1281 429 -881
<< ndiff >>
rect -487 1331 -429 1343
rect -487 955 -475 1331
rect -441 955 -429 1331
rect -487 943 -429 955
rect -29 1331 29 1343
rect -29 955 -17 1331
rect 17 955 29 1331
rect -29 943 29 955
rect 429 1331 487 1343
rect 429 955 441 1331
rect 475 955 487 1331
rect 429 943 487 955
rect -487 775 -429 787
rect -487 399 -475 775
rect -441 399 -429 775
rect -487 387 -429 399
rect -29 775 29 787
rect -29 399 -17 775
rect 17 399 29 775
rect -29 387 29 399
rect 429 775 487 787
rect 429 399 441 775
rect 475 399 487 775
rect 429 387 487 399
rect -487 219 -429 231
rect -487 -157 -475 219
rect -441 -157 -429 219
rect -487 -169 -429 -157
rect -29 219 29 231
rect -29 -157 -17 219
rect 17 -157 29 219
rect -29 -169 29 -157
rect 429 219 487 231
rect 429 -157 441 219
rect 475 -157 487 219
rect 429 -169 487 -157
rect -487 -337 -429 -325
rect -487 -713 -475 -337
rect -441 -713 -429 -337
rect -487 -725 -429 -713
rect -29 -337 29 -325
rect -29 -713 -17 -337
rect 17 -713 29 -337
rect -29 -725 29 -713
rect 429 -337 487 -325
rect 429 -713 441 -337
rect 475 -713 487 -337
rect 429 -725 487 -713
rect -487 -893 -429 -881
rect -487 -1269 -475 -893
rect -441 -1269 -429 -893
rect -487 -1281 -429 -1269
rect -29 -893 29 -881
rect -29 -1269 -17 -893
rect 17 -1269 29 -893
rect -29 -1281 29 -1269
rect 429 -893 487 -881
rect 429 -1269 441 -893
rect 475 -1269 487 -893
rect 429 -1281 487 -1269
<< ndiffc >>
rect -475 955 -441 1331
rect -17 955 17 1331
rect 441 955 475 1331
rect -475 399 -441 775
rect -17 399 17 775
rect 441 399 475 775
rect -475 -157 -441 219
rect -17 -157 17 219
rect 441 -157 475 219
rect -475 -713 -441 -337
rect -17 -713 17 -337
rect 441 -713 475 -337
rect -475 -1269 -441 -893
rect -17 -1269 17 -893
rect 441 -1269 475 -893
<< psubdiff >>
rect -589 1421 -493 1455
rect 493 1421 589 1455
rect -589 1359 -555 1421
rect 555 1359 589 1421
rect -589 -1421 -555 -1359
rect 555 -1421 589 -1359
rect -589 -1455 -493 -1421
rect 493 -1455 589 -1421
<< psubdiffcont >>
rect -493 1421 493 1455
rect -589 -1359 -555 1359
rect 555 -1359 589 1359
rect -493 -1455 493 -1421
<< poly >>
rect -429 1343 -29 1369
rect 29 1343 429 1369
rect -429 905 -29 943
rect -429 871 -413 905
rect -45 871 -29 905
rect -429 855 -29 871
rect 29 905 429 943
rect 29 871 45 905
rect 413 871 429 905
rect 29 855 429 871
rect -429 787 -29 813
rect 29 787 429 813
rect -429 349 -29 387
rect -429 315 -413 349
rect -45 315 -29 349
rect -429 299 -29 315
rect 29 349 429 387
rect 29 315 45 349
rect 413 315 429 349
rect 29 299 429 315
rect -429 231 -29 257
rect 29 231 429 257
rect -429 -207 -29 -169
rect -429 -241 -413 -207
rect -45 -241 -29 -207
rect -429 -257 -29 -241
rect 29 -207 429 -169
rect 29 -241 45 -207
rect 413 -241 429 -207
rect 29 -257 429 -241
rect -429 -325 -29 -299
rect 29 -325 429 -299
rect -429 -763 -29 -725
rect -429 -797 -413 -763
rect -45 -797 -29 -763
rect -429 -813 -29 -797
rect 29 -763 429 -725
rect 29 -797 45 -763
rect 413 -797 429 -763
rect 29 -813 429 -797
rect -429 -881 -29 -855
rect 29 -881 429 -855
rect -429 -1319 -29 -1281
rect -429 -1353 -413 -1319
rect -45 -1353 -29 -1319
rect -429 -1369 -29 -1353
rect 29 -1319 429 -1281
rect 29 -1353 45 -1319
rect 413 -1353 429 -1319
rect 29 -1369 429 -1353
<< polycont >>
rect -413 871 -45 905
rect 45 871 413 905
rect -413 315 -45 349
rect 45 315 413 349
rect -413 -241 -45 -207
rect 45 -241 413 -207
rect -413 -797 -45 -763
rect 45 -797 413 -763
rect -413 -1353 -45 -1319
rect 45 -1353 413 -1319
<< locali >>
rect -589 1421 -493 1455
rect 493 1421 589 1455
rect -589 1359 -555 1421
rect 555 1359 589 1421
rect -475 1331 -441 1347
rect -475 939 -441 955
rect -17 1331 17 1347
rect -17 939 17 955
rect 441 1331 475 1347
rect 441 939 475 955
rect -429 871 -413 905
rect -45 871 -29 905
rect 29 871 45 905
rect 413 871 429 905
rect -475 775 -441 791
rect -475 383 -441 399
rect -17 775 17 791
rect -17 383 17 399
rect 441 775 475 791
rect 441 383 475 399
rect -429 315 -413 349
rect -45 315 -29 349
rect 29 315 45 349
rect 413 315 429 349
rect -475 219 -441 235
rect -475 -173 -441 -157
rect -17 219 17 235
rect -17 -173 17 -157
rect 441 219 475 235
rect 441 -173 475 -157
rect -429 -241 -413 -207
rect -45 -241 -29 -207
rect 29 -241 45 -207
rect 413 -241 429 -207
rect -475 -337 -441 -321
rect -475 -729 -441 -713
rect -17 -337 17 -321
rect -17 -729 17 -713
rect 441 -337 475 -321
rect 441 -729 475 -713
rect -429 -797 -413 -763
rect -45 -797 -29 -763
rect 29 -797 45 -763
rect 413 -797 429 -763
rect -475 -893 -441 -877
rect -475 -1285 -441 -1269
rect -17 -893 17 -877
rect -17 -1285 17 -1269
rect 441 -893 475 -877
rect 441 -1285 475 -1269
rect -429 -1353 -413 -1319
rect -45 -1353 -29 -1319
rect 29 -1353 45 -1319
rect 413 -1353 429 -1319
rect -589 -1421 -555 -1359
rect 555 -1421 589 -1359
rect -589 -1455 -493 -1421
rect 493 -1455 589 -1421
<< viali >>
rect -475 955 -441 1331
rect -17 955 17 1331
rect 441 955 475 1331
rect -413 871 -45 905
rect 45 871 413 905
rect -475 399 -441 775
rect -17 399 17 775
rect 441 399 475 775
rect -413 315 -45 349
rect 45 315 413 349
rect -475 -157 -441 219
rect -17 -157 17 219
rect 441 -157 475 219
rect -413 -241 -45 -207
rect 45 -241 413 -207
rect -475 -713 -441 -337
rect -17 -713 17 -337
rect 441 -713 475 -337
rect -413 -797 -45 -763
rect 45 -797 413 -763
rect -475 -1269 -441 -893
rect -17 -1269 17 -893
rect 441 -1269 475 -893
rect -413 -1353 -45 -1319
rect 45 -1353 413 -1319
<< metal1 >>
rect -481 1331 -435 1343
rect -481 955 -475 1331
rect -441 955 -435 1331
rect -481 943 -435 955
rect -23 1331 23 1343
rect -23 955 -17 1331
rect 17 955 23 1331
rect -23 943 23 955
rect 435 1331 481 1343
rect 435 955 441 1331
rect 475 955 481 1331
rect 435 943 481 955
rect -425 905 -33 911
rect -425 871 -413 905
rect -45 871 -33 905
rect -425 865 -33 871
rect 33 905 425 911
rect 33 871 45 905
rect 413 871 425 905
rect 33 865 425 871
rect -481 775 -435 787
rect -481 399 -475 775
rect -441 399 -435 775
rect -481 387 -435 399
rect -23 775 23 787
rect -23 399 -17 775
rect 17 399 23 775
rect -23 387 23 399
rect 435 775 481 787
rect 435 399 441 775
rect 475 399 481 775
rect 435 387 481 399
rect -425 349 -33 355
rect -425 315 -413 349
rect -45 315 -33 349
rect -425 309 -33 315
rect 33 349 425 355
rect 33 315 45 349
rect 413 315 425 349
rect 33 309 425 315
rect -481 219 -435 231
rect -481 -157 -475 219
rect -441 -157 -435 219
rect -481 -169 -435 -157
rect -23 219 23 231
rect -23 -157 -17 219
rect 17 -157 23 219
rect -23 -169 23 -157
rect 435 219 481 231
rect 435 -157 441 219
rect 475 -157 481 219
rect 435 -169 481 -157
rect -425 -207 -33 -201
rect -425 -241 -413 -207
rect -45 -241 -33 -207
rect -425 -247 -33 -241
rect 33 -207 425 -201
rect 33 -241 45 -207
rect 413 -241 425 -207
rect 33 -247 425 -241
rect -481 -337 -435 -325
rect -481 -713 -475 -337
rect -441 -713 -435 -337
rect -481 -725 -435 -713
rect -23 -337 23 -325
rect -23 -713 -17 -337
rect 17 -713 23 -337
rect -23 -725 23 -713
rect 435 -337 481 -325
rect 435 -713 441 -337
rect 475 -713 481 -337
rect 435 -725 481 -713
rect -425 -763 -33 -757
rect -425 -797 -413 -763
rect -45 -797 -33 -763
rect -425 -803 -33 -797
rect 33 -763 425 -757
rect 33 -797 45 -763
rect 413 -797 425 -763
rect 33 -803 425 -797
rect -481 -893 -435 -881
rect -481 -1269 -475 -893
rect -441 -1269 -435 -893
rect -481 -1281 -435 -1269
rect -23 -893 23 -881
rect -23 -1269 -17 -893
rect 17 -1269 23 -893
rect -23 -1281 23 -1269
rect 435 -893 481 -881
rect 435 -1269 441 -893
rect 475 -1269 481 -893
rect 435 -1281 481 -1269
rect -425 -1319 -33 -1313
rect -425 -1353 -413 -1319
rect -45 -1353 -33 -1319
rect -425 -1359 -33 -1353
rect 33 -1319 425 -1313
rect 33 -1353 45 -1319
rect 413 -1353 425 -1319
rect 33 -1359 425 -1353
<< properties >>
string FIXED_BBOX -572 -1438 572 1438
string gencell sky130_fd_pr__nfet_01v8_lvt
string library sky130
string parameters w 2 l 2 m 5 nf 2 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 0 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
