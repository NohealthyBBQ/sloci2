magic
tech sky130A
magscale 1 2
timestamp 1662511141
<< locali >>
rect 520 1220 580 1300
<< metal1 >>
rect 50 1060 60 1120
rect 140 1060 150 1120
rect 550 1060 560 1120
rect 640 1060 650 1120
rect 1070 1060 1080 1120
rect 1160 1060 1170 1120
rect 290 740 300 800
rect 380 740 390 800
rect 810 740 820 800
rect 900 740 910 800
rect 320 664 400 698
rect 50 500 60 560
rect 140 500 150 560
rect 310 180 320 240
rect 400 180 410 240
rect 318 108 398 142
rect 440 100 500 700
rect 570 666 650 700
rect 834 666 914 700
rect 570 500 580 560
rect 660 500 670 560
rect 1090 520 1100 580
rect 1180 520 1190 580
rect 810 180 820 240
rect 900 180 910 240
rect 574 112 654 146
rect 830 108 910 142
<< via1 >>
rect 60 1060 140 1120
rect 560 1060 640 1120
rect 1080 1060 1160 1120
rect 300 740 380 800
rect 820 740 900 800
rect 60 500 140 560
rect 320 180 400 240
rect 580 500 660 560
rect 1100 520 1180 580
rect 820 180 900 240
<< metal2 >>
rect -100 1120 1160 1140
rect -100 1060 60 1120
rect 140 1060 560 1120
rect 640 1060 1080 1120
rect -100 1040 1160 1060
rect -100 580 -60 1040
rect 300 800 380 810
rect 820 800 900 810
rect 1300 800 1340 820
rect 280 740 300 800
rect 380 740 820 800
rect 900 740 1360 800
rect 300 730 380 740
rect 820 730 1360 740
rect 880 720 1360 730
rect 1100 580 1180 590
rect -100 560 1100 580
rect -100 500 60 560
rect 140 500 580 560
rect 660 520 1100 560
rect 660 500 1180 520
rect -100 490 140 500
rect 580 490 660 500
rect -100 480 80 490
rect 300 240 900 260
rect 1300 240 1340 720
rect 300 180 320 240
rect 400 180 820 240
rect 900 180 1360 240
rect 300 160 1360 180
use sky130_fd_pr__nfet_01v8_lvt_T7FZYG  sky130_fd_pr__nfet_01v8_lvt_T7FZYG_0
timestamp 1662510765
transform 1 0 614 0 1 628
box -683 -657 683 657
<< labels >>
rlabel metal2 900 720 1360 800 3 D
rlabel metal2 -100 480 -60 1140 7 S
rlabel space 440 100 500 705 0 G
rlabel locali 520 1220 580 1300 1 B
<< end >>
