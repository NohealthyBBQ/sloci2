magic
tech sky130A
magscale 1 2
timestamp 1662510765
<< pwell >>
rect -683 -657 683 657
<< nmoslvt >>
rect -487 109 -287 509
rect -229 109 -29 509
rect 29 109 229 509
rect 287 109 487 509
rect -487 -447 -287 -47
rect -229 -447 -29 -47
rect 29 -447 229 -47
rect 287 -447 487 -47
<< ndiff >>
rect -545 497 -487 509
rect -545 121 -533 497
rect -499 121 -487 497
rect -545 109 -487 121
rect -287 497 -229 509
rect -287 121 -275 497
rect -241 121 -229 497
rect -287 109 -229 121
rect -29 497 29 509
rect -29 121 -17 497
rect 17 121 29 497
rect -29 109 29 121
rect 229 497 287 509
rect 229 121 241 497
rect 275 121 287 497
rect 229 109 287 121
rect 487 497 545 509
rect 487 121 499 497
rect 533 121 545 497
rect 487 109 545 121
rect -545 -59 -487 -47
rect -545 -435 -533 -59
rect -499 -435 -487 -59
rect -545 -447 -487 -435
rect -287 -59 -229 -47
rect -287 -435 -275 -59
rect -241 -435 -229 -59
rect -287 -447 -229 -435
rect -29 -59 29 -47
rect -29 -435 -17 -59
rect 17 -435 29 -59
rect -29 -447 29 -435
rect 229 -59 287 -47
rect 229 -435 241 -59
rect 275 -435 287 -59
rect 229 -447 287 -435
rect 487 -59 545 -47
rect 487 -435 499 -59
rect 533 -435 545 -59
rect 487 -447 545 -435
<< ndiffc >>
rect -533 121 -499 497
rect -275 121 -241 497
rect -17 121 17 497
rect 241 121 275 497
rect 499 121 533 497
rect -533 -435 -499 -59
rect -275 -435 -241 -59
rect -17 -435 17 -59
rect 241 -435 275 -59
rect 499 -435 533 -59
<< psubdiff >>
rect -647 587 -551 621
rect 551 587 647 621
rect -647 525 -613 587
rect 613 525 647 587
rect -647 -587 -613 -525
rect 613 -587 647 -525
rect -647 -621 -551 -587
rect 551 -621 647 -587
<< psubdiffcont >>
rect -551 587 551 621
rect -647 -525 -613 525
rect 613 -525 647 525
rect -551 -621 551 -587
<< poly >>
rect -487 509 -287 535
rect -229 509 -29 535
rect 29 509 229 535
rect 287 509 487 535
rect -487 71 -287 109
rect -487 37 -471 71
rect -303 37 -287 71
rect -487 21 -287 37
rect -229 71 -29 109
rect -229 37 -213 71
rect -45 37 -29 71
rect -229 21 -29 37
rect 29 71 229 109
rect 29 37 45 71
rect 213 37 229 71
rect 29 21 229 37
rect 287 71 487 109
rect 287 37 303 71
rect 471 37 487 71
rect 287 21 487 37
rect -487 -47 -287 -21
rect -229 -47 -29 -21
rect 29 -47 229 -21
rect 287 -47 487 -21
rect -487 -485 -287 -447
rect -487 -519 -471 -485
rect -303 -519 -287 -485
rect -487 -535 -287 -519
rect -229 -485 -29 -447
rect -229 -519 -213 -485
rect -45 -519 -29 -485
rect -229 -535 -29 -519
rect 29 -485 229 -447
rect 29 -519 45 -485
rect 213 -519 229 -485
rect 29 -535 229 -519
rect 287 -485 487 -447
rect 287 -519 303 -485
rect 471 -519 487 -485
rect 287 -535 487 -519
<< polycont >>
rect -471 37 -303 71
rect -213 37 -45 71
rect 45 37 213 71
rect 303 37 471 71
rect -471 -519 -303 -485
rect -213 -519 -45 -485
rect 45 -519 213 -485
rect 303 -519 471 -485
<< locali >>
rect -647 587 -551 621
rect 551 587 647 621
rect -647 525 -613 587
rect 613 525 647 587
rect -533 497 -499 513
rect -533 105 -499 121
rect -275 497 -241 513
rect -275 105 -241 121
rect -17 497 17 513
rect -17 105 17 121
rect 241 497 275 513
rect 241 105 275 121
rect 499 497 533 513
rect 499 105 533 121
rect -487 37 -471 71
rect -303 37 -287 71
rect -229 37 -213 71
rect -45 37 -29 71
rect 29 37 45 71
rect 213 37 229 71
rect 287 37 303 71
rect 471 37 487 71
rect -533 -59 -499 -43
rect -533 -451 -499 -435
rect -275 -59 -241 -43
rect -275 -451 -241 -435
rect -17 -59 17 -43
rect -17 -451 17 -435
rect 241 -59 275 -43
rect 241 -451 275 -435
rect 499 -59 533 -43
rect 499 -451 533 -435
rect -487 -519 -471 -485
rect -303 -519 -287 -485
rect -229 -519 -213 -485
rect -45 -519 -29 -485
rect 29 -519 45 -485
rect 213 -519 229 -485
rect 287 -519 303 -485
rect 471 -519 487 -485
rect -647 -587 -613 -525
rect 613 -587 647 -525
rect -647 -621 -551 -587
rect 551 -621 647 -587
<< viali >>
rect -533 121 -499 497
rect -275 121 -241 497
rect -17 121 17 497
rect 241 121 275 497
rect 499 121 533 497
rect -471 37 -303 71
rect -213 37 -45 71
rect 45 37 213 71
rect 303 37 471 71
rect -533 -435 -499 -59
rect -275 -435 -241 -59
rect -17 -435 17 -59
rect 241 -435 275 -59
rect 499 -435 533 -59
rect -471 -519 -303 -485
rect -213 -519 -45 -485
rect 45 -519 213 -485
rect 303 -519 471 -485
<< metal1 >>
rect -539 497 -493 509
rect -539 121 -533 497
rect -499 121 -493 497
rect -539 109 -493 121
rect -281 497 -235 509
rect -281 121 -275 497
rect -241 121 -235 497
rect -281 109 -235 121
rect -23 497 23 509
rect -23 121 -17 497
rect 17 121 23 497
rect -23 109 23 121
rect 235 497 281 509
rect 235 121 241 497
rect 275 121 281 497
rect 235 109 281 121
rect 493 497 539 509
rect 493 121 499 497
rect 533 121 539 497
rect 493 109 539 121
rect -483 71 -291 77
rect -483 37 -471 71
rect -303 37 -291 71
rect -483 31 -291 37
rect -225 71 -33 77
rect -225 37 -213 71
rect -45 37 -33 71
rect -225 31 -33 37
rect 33 71 225 77
rect 33 37 45 71
rect 213 37 225 71
rect 33 31 225 37
rect 291 71 483 77
rect 291 37 303 71
rect 471 37 483 71
rect 291 31 483 37
rect -539 -59 -493 -47
rect -539 -435 -533 -59
rect -499 -435 -493 -59
rect -539 -447 -493 -435
rect -281 -59 -235 -47
rect -281 -435 -275 -59
rect -241 -435 -235 -59
rect -281 -447 -235 -435
rect -23 -59 23 -47
rect -23 -435 -17 -59
rect 17 -435 23 -59
rect -23 -447 23 -435
rect 235 -59 281 -47
rect 235 -435 241 -59
rect 275 -435 281 -59
rect 235 -447 281 -435
rect 493 -59 539 -47
rect 493 -435 499 -59
rect 533 -435 539 -59
rect 493 -447 539 -435
rect -483 -485 -291 -479
rect -483 -519 -471 -485
rect -303 -519 -291 -485
rect -483 -525 -291 -519
rect -225 -485 -33 -479
rect -225 -519 -213 -485
rect -45 -519 -33 -485
rect -225 -525 -33 -519
rect 33 -485 225 -479
rect 33 -519 45 -485
rect 213 -519 225 -485
rect 33 -525 225 -519
rect 291 -485 483 -479
rect 291 -519 303 -485
rect 471 -519 483 -485
rect 291 -525 483 -519
<< properties >>
string FIXED_BBOX -630 -604 630 604
string gencell sky130_fd_pr__nfet_01v8_lvt
string library sky130
string parameters w 2 l 1 m 2 nf 4 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 0 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
