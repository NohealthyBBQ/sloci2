magic
tech sky130A
magscale 1 2
timestamp 1661909182
<< nwell >>
rect -2129 -298 2129 264
<< pmoslvt >>
rect -2035 -236 -1835 164
rect -1777 -236 -1577 164
rect -1519 -236 -1319 164
rect -1261 -236 -1061 164
rect -1003 -236 -803 164
rect -745 -236 -545 164
rect -487 -236 -287 164
rect -229 -236 -29 164
rect 29 -236 229 164
rect 287 -236 487 164
rect 545 -236 745 164
rect 803 -236 1003 164
rect 1061 -236 1261 164
rect 1319 -236 1519 164
rect 1577 -236 1777 164
rect 1835 -236 2035 164
<< pdiff >>
rect -2093 152 -2035 164
rect -2093 -224 -2081 152
rect -2047 -224 -2035 152
rect -2093 -236 -2035 -224
rect -1835 152 -1777 164
rect -1835 -224 -1823 152
rect -1789 -224 -1777 152
rect -1835 -236 -1777 -224
rect -1577 152 -1519 164
rect -1577 -224 -1565 152
rect -1531 -224 -1519 152
rect -1577 -236 -1519 -224
rect -1319 152 -1261 164
rect -1319 -224 -1307 152
rect -1273 -224 -1261 152
rect -1319 -236 -1261 -224
rect -1061 152 -1003 164
rect -1061 -224 -1049 152
rect -1015 -224 -1003 152
rect -1061 -236 -1003 -224
rect -803 152 -745 164
rect -803 -224 -791 152
rect -757 -224 -745 152
rect -803 -236 -745 -224
rect -545 152 -487 164
rect -545 -224 -533 152
rect -499 -224 -487 152
rect -545 -236 -487 -224
rect -287 152 -229 164
rect -287 -224 -275 152
rect -241 -224 -229 152
rect -287 -236 -229 -224
rect -29 152 29 164
rect -29 -224 -17 152
rect 17 -224 29 152
rect -29 -236 29 -224
rect 229 152 287 164
rect 229 -224 241 152
rect 275 -224 287 152
rect 229 -236 287 -224
rect 487 152 545 164
rect 487 -224 499 152
rect 533 -224 545 152
rect 487 -236 545 -224
rect 745 152 803 164
rect 745 -224 757 152
rect 791 -224 803 152
rect 745 -236 803 -224
rect 1003 152 1061 164
rect 1003 -224 1015 152
rect 1049 -224 1061 152
rect 1003 -236 1061 -224
rect 1261 152 1319 164
rect 1261 -224 1273 152
rect 1307 -224 1319 152
rect 1261 -236 1319 -224
rect 1519 152 1577 164
rect 1519 -224 1531 152
rect 1565 -224 1577 152
rect 1519 -236 1577 -224
rect 1777 152 1835 164
rect 1777 -224 1789 152
rect 1823 -224 1835 152
rect 1777 -236 1835 -224
rect 2035 152 2093 164
rect 2035 -224 2047 152
rect 2081 -224 2093 152
rect 2035 -236 2093 -224
<< pdiffc >>
rect -2081 -224 -2047 152
rect -1823 -224 -1789 152
rect -1565 -224 -1531 152
rect -1307 -224 -1273 152
rect -1049 -224 -1015 152
rect -791 -224 -757 152
rect -533 -224 -499 152
rect -275 -224 -241 152
rect -17 -224 17 152
rect 241 -224 275 152
rect 499 -224 533 152
rect 757 -224 791 152
rect 1015 -224 1049 152
rect 1273 -224 1307 152
rect 1531 -224 1565 152
rect 1789 -224 1823 152
rect 2047 -224 2081 152
<< poly >>
rect -2035 245 -1835 261
rect -2035 211 -2019 245
rect -1851 211 -1835 245
rect -2035 164 -1835 211
rect -1777 245 -1577 261
rect -1777 211 -1761 245
rect -1593 211 -1577 245
rect -1777 164 -1577 211
rect -1519 245 -1319 261
rect -1519 211 -1503 245
rect -1335 211 -1319 245
rect -1519 164 -1319 211
rect -1261 245 -1061 261
rect -1261 211 -1245 245
rect -1077 211 -1061 245
rect -1261 164 -1061 211
rect -1003 245 -803 261
rect -1003 211 -987 245
rect -819 211 -803 245
rect -1003 164 -803 211
rect -745 245 -545 261
rect -745 211 -729 245
rect -561 211 -545 245
rect -745 164 -545 211
rect -487 245 -287 261
rect -487 211 -471 245
rect -303 211 -287 245
rect -487 164 -287 211
rect -229 245 -29 261
rect -229 211 -213 245
rect -45 211 -29 245
rect -229 164 -29 211
rect 29 245 229 261
rect 29 211 45 245
rect 213 211 229 245
rect 29 164 229 211
rect 287 245 487 261
rect 287 211 303 245
rect 471 211 487 245
rect 287 164 487 211
rect 545 245 745 261
rect 545 211 561 245
rect 729 211 745 245
rect 545 164 745 211
rect 803 245 1003 261
rect 803 211 819 245
rect 987 211 1003 245
rect 803 164 1003 211
rect 1061 245 1261 261
rect 1061 211 1077 245
rect 1245 211 1261 245
rect 1061 164 1261 211
rect 1319 245 1519 261
rect 1319 211 1335 245
rect 1503 211 1519 245
rect 1319 164 1519 211
rect 1577 245 1777 261
rect 1577 211 1593 245
rect 1761 211 1777 245
rect 1577 164 1777 211
rect 1835 245 2035 261
rect 1835 211 1851 245
rect 2019 211 2035 245
rect 1835 164 2035 211
rect -2035 -262 -1835 -236
rect -1777 -262 -1577 -236
rect -1519 -262 -1319 -236
rect -1261 -262 -1061 -236
rect -1003 -262 -803 -236
rect -745 -262 -545 -236
rect -487 -262 -287 -236
rect -229 -262 -29 -236
rect 29 -262 229 -236
rect 287 -262 487 -236
rect 545 -262 745 -236
rect 803 -262 1003 -236
rect 1061 -262 1261 -236
rect 1319 -262 1519 -236
rect 1577 -262 1777 -236
rect 1835 -262 2035 -236
<< polycont >>
rect -2019 211 -1851 245
rect -1761 211 -1593 245
rect -1503 211 -1335 245
rect -1245 211 -1077 245
rect -987 211 -819 245
rect -729 211 -561 245
rect -471 211 -303 245
rect -213 211 -45 245
rect 45 211 213 245
rect 303 211 471 245
rect 561 211 729 245
rect 819 211 987 245
rect 1077 211 1245 245
rect 1335 211 1503 245
rect 1593 211 1761 245
rect 1851 211 2019 245
<< locali >>
rect -2035 211 -2019 245
rect -1851 211 -1835 245
rect -1777 211 -1761 245
rect -1593 211 -1577 245
rect -1519 211 -1503 245
rect -1335 211 -1319 245
rect -1261 211 -1245 245
rect -1077 211 -1061 245
rect -1003 211 -987 245
rect -819 211 -803 245
rect -745 211 -729 245
rect -561 211 -545 245
rect -487 211 -471 245
rect -303 211 -287 245
rect -229 211 -213 245
rect -45 211 -29 245
rect 29 211 45 245
rect 213 211 229 245
rect 287 211 303 245
rect 471 211 487 245
rect 545 211 561 245
rect 729 211 745 245
rect 803 211 819 245
rect 987 211 1003 245
rect 1061 211 1077 245
rect 1245 211 1261 245
rect 1319 211 1335 245
rect 1503 211 1519 245
rect 1577 211 1593 245
rect 1761 211 1777 245
rect 1835 211 1851 245
rect 2019 211 2035 245
rect -2081 152 -2047 168
rect -2081 -240 -2047 -224
rect -1823 152 -1789 168
rect -1823 -240 -1789 -224
rect -1565 152 -1531 168
rect -1565 -240 -1531 -224
rect -1307 152 -1273 168
rect -1307 -240 -1273 -224
rect -1049 152 -1015 168
rect -1049 -240 -1015 -224
rect -791 152 -757 168
rect -791 -240 -757 -224
rect -533 152 -499 168
rect -533 -240 -499 -224
rect -275 152 -241 168
rect -275 -240 -241 -224
rect -17 152 17 168
rect -17 -240 17 -224
rect 241 152 275 168
rect 241 -240 275 -224
rect 499 152 533 168
rect 499 -240 533 -224
rect 757 152 791 168
rect 757 -240 791 -224
rect 1015 152 1049 168
rect 1015 -240 1049 -224
rect 1273 152 1307 168
rect 1273 -240 1307 -224
rect 1531 152 1565 168
rect 1531 -240 1565 -224
rect 1789 152 1823 168
rect 1789 -240 1823 -224
rect 2047 152 2081 168
rect 2047 -240 2081 -224
<< viali >>
rect -2019 211 -1851 245
rect -1761 211 -1593 245
rect -1503 211 -1335 245
rect -1245 211 -1077 245
rect -987 211 -819 245
rect -729 211 -561 245
rect -471 211 -303 245
rect -213 211 -45 245
rect 45 211 213 245
rect 303 211 471 245
rect 561 211 729 245
rect 819 211 987 245
rect 1077 211 1245 245
rect 1335 211 1503 245
rect 1593 211 1761 245
rect 1851 211 2019 245
rect -2081 -224 -2047 152
rect -1823 -224 -1789 152
rect -1565 -224 -1531 152
rect -1307 -224 -1273 152
rect -1049 -224 -1015 152
rect -791 -224 -757 152
rect -533 -224 -499 152
rect -275 -224 -241 152
rect -17 -224 17 152
rect 241 -224 275 152
rect 499 -224 533 152
rect 757 -224 791 152
rect 1015 -224 1049 152
rect 1273 -224 1307 152
rect 1531 -224 1565 152
rect 1789 -224 1823 152
rect 2047 -224 2081 152
<< metal1 >>
rect -2031 245 -1839 251
rect -2031 211 -2019 245
rect -1851 211 -1839 245
rect -2031 205 -1839 211
rect -1773 245 -1581 251
rect -1773 211 -1761 245
rect -1593 211 -1581 245
rect -1773 205 -1581 211
rect -1515 245 -1323 251
rect -1515 211 -1503 245
rect -1335 211 -1323 245
rect -1515 205 -1323 211
rect -1257 245 -1065 251
rect -1257 211 -1245 245
rect -1077 211 -1065 245
rect -1257 205 -1065 211
rect -999 245 -807 251
rect -999 211 -987 245
rect -819 211 -807 245
rect -999 205 -807 211
rect -741 245 -549 251
rect -741 211 -729 245
rect -561 211 -549 245
rect -741 205 -549 211
rect -483 245 -291 251
rect -483 211 -471 245
rect -303 211 -291 245
rect -483 205 -291 211
rect -225 245 -33 251
rect -225 211 -213 245
rect -45 211 -33 245
rect -225 205 -33 211
rect 33 245 225 251
rect 33 211 45 245
rect 213 211 225 245
rect 33 205 225 211
rect 291 245 483 251
rect 291 211 303 245
rect 471 211 483 245
rect 291 205 483 211
rect 549 245 741 251
rect 549 211 561 245
rect 729 211 741 245
rect 549 205 741 211
rect 807 245 999 251
rect 807 211 819 245
rect 987 211 999 245
rect 807 205 999 211
rect 1065 245 1257 251
rect 1065 211 1077 245
rect 1245 211 1257 245
rect 1065 205 1257 211
rect 1323 245 1515 251
rect 1323 211 1335 245
rect 1503 211 1515 245
rect 1323 205 1515 211
rect 1581 245 1773 251
rect 1581 211 1593 245
rect 1761 211 1773 245
rect 1581 205 1773 211
rect 1839 245 2031 251
rect 1839 211 1851 245
rect 2019 211 2031 245
rect 1839 205 2031 211
rect -2087 152 -2041 164
rect -2087 -224 -2081 152
rect -2047 -224 -2041 152
rect -2087 -236 -2041 -224
rect -1829 152 -1783 164
rect -1829 -224 -1823 152
rect -1789 -224 -1783 152
rect -1829 -236 -1783 -224
rect -1571 152 -1525 164
rect -1571 -224 -1565 152
rect -1531 -224 -1525 152
rect -1571 -236 -1525 -224
rect -1313 152 -1267 164
rect -1313 -224 -1307 152
rect -1273 -224 -1267 152
rect -1313 -236 -1267 -224
rect -1055 152 -1009 164
rect -1055 -224 -1049 152
rect -1015 -224 -1009 152
rect -1055 -236 -1009 -224
rect -797 152 -751 164
rect -797 -224 -791 152
rect -757 -224 -751 152
rect -797 -236 -751 -224
rect -539 152 -493 164
rect -539 -224 -533 152
rect -499 -224 -493 152
rect -539 -236 -493 -224
rect -281 152 -235 164
rect -281 -224 -275 152
rect -241 -224 -235 152
rect -281 -236 -235 -224
rect -23 152 23 164
rect -23 -224 -17 152
rect 17 -224 23 152
rect -23 -236 23 -224
rect 235 152 281 164
rect 235 -224 241 152
rect 275 -224 281 152
rect 235 -236 281 -224
rect 493 152 539 164
rect 493 -224 499 152
rect 533 -224 539 152
rect 493 -236 539 -224
rect 751 152 797 164
rect 751 -224 757 152
rect 791 -224 797 152
rect 751 -236 797 -224
rect 1009 152 1055 164
rect 1009 -224 1015 152
rect 1049 -224 1055 152
rect 1009 -236 1055 -224
rect 1267 152 1313 164
rect 1267 -224 1273 152
rect 1307 -224 1313 152
rect 1267 -236 1313 -224
rect 1525 152 1571 164
rect 1525 -224 1531 152
rect 1565 -224 1571 152
rect 1525 -236 1571 -224
rect 1783 152 1829 164
rect 1783 -224 1789 152
rect 1823 -224 1829 152
rect 1783 -236 1829 -224
rect 2041 152 2087 164
rect 2041 -224 2047 152
rect 2081 -224 2087 152
rect 2041 -236 2087 -224
<< properties >>
string gencell sky130_fd_pr__pfet_01v8_lvt
string library sky130
string parameters w 2 l 1 m 1 nf 16 diffcov 100 polycov 100 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 0 poverlap 0 doverlap 1 lmin 0.35 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
