magic
tech sky130A
magscale 1 2
timestamp 1672329920
<< locali >>
rect 14600 3780 15000 3800
rect 14600 3320 14620 3780
rect 14980 3320 15000 3780
rect 14600 3300 15000 3320
rect 25300 2040 25860 3320
<< viali >>
rect 14620 3320 14980 3780
<< metal1 >>
rect 14614 3780 14986 3792
rect 14610 3320 14620 3780
rect 14980 3320 14990 3780
rect 14614 3308 14986 3320
rect 15000 1400 15200 2400
rect 25400 400 25600 1400
rect 15000 -1000 15200 0
rect 25400 -2200 25600 -1200
rect 15000 -3400 15200 -2400
rect 25400 -4800 25600 -3800
rect 15000 -6000 15200 -5000
rect 25400 -7200 25600 -6200
rect 15000 -8400 15200 -7400
rect 25400 -9600 25600 -8600
rect 15000 -11000 15200 -10000
rect 25400 -12200 25600 -11200
rect 14840 -13120 14940 -12720
rect 15830 -13260 15840 -13180
rect 15920 -13260 15930 -13180
rect 14820 -13900 14860 -13420
rect 16920 -13540 16960 -13060
rect 15830 -13620 15840 -13540
rect 15920 -13620 15930 -13540
rect 15830 -13980 15840 -13900
rect 15920 -13980 15930 -13900
rect 14820 -14620 14860 -14140
rect 16920 -14260 16960 -13780
rect 15830 -14340 15840 -14260
rect 15920 -14340 15930 -14260
rect 15830 -14700 15840 -14620
rect 15920 -14700 15930 -14620
rect 14820 -15340 14860 -14860
rect 16920 -14980 16960 -14500
rect 15830 -15060 15840 -14980
rect 15920 -15060 15930 -14980
rect 15830 -15420 15840 -15340
rect 15920 -15420 15930 -15340
rect 14820 -16220 15000 -15580
rect 16920 -15680 16960 -15220
rect 15830 -15780 15840 -15700
rect 15920 -15780 15930 -15700
rect 14820 -16380 14840 -16220
rect 14980 -16380 15000 -16220
<< via1 >>
rect 14620 3320 14980 3780
rect 15840 -13260 15920 -13180
rect 15840 -13620 15920 -13540
rect 15840 -13980 15920 -13900
rect 15840 -14340 15920 -14260
rect 15840 -14700 15920 -14620
rect 15840 -15060 15920 -14980
rect 15840 -15420 15920 -15340
rect 15840 -15780 15920 -15700
rect 14840 -16380 14980 -16220
<< metal2 >>
rect 14620 3780 14980 3790
rect 14620 3310 14980 3320
rect 15840 -13180 15920 -13160
rect 15840 -13540 15920 -13260
rect 15840 -13900 15920 -13620
rect 15840 -14260 15920 -13980
rect 15840 -14620 15920 -14340
rect 15840 -14980 15920 -14700
rect 15840 -15340 15920 -15060
rect 15840 -15700 15920 -15420
rect 15840 -15800 15920 -15780
rect 14840 -16220 14980 -16210
rect 14840 -16390 14980 -16380
<< via2 >>
rect 14620 3320 14980 3780
rect 14840 -16380 14980 -16220
<< metal3 >>
rect 6800 5600 9000 6200
rect 14000 3780 15000 3800
rect 14000 3400 14620 3780
rect 14600 3320 14620 3400
rect 14980 3320 15000 3780
rect 14600 3300 15000 3320
rect 7000 -13400 8600 -12800
rect 14830 -16220 14990 -16215
rect 14830 -16380 14840 -16220
rect 14980 -16380 14990 -16220
rect 14830 -16385 14990 -16380
<< via3 >>
rect 14840 -16380 14980 -16220
<< metal4 >>
rect 6400 -16200 6600 -15400
rect 13200 -16200 13400 -15400
rect 6400 -16220 15000 -16200
rect 6400 -16380 14840 -16220
rect 14980 -16380 15000 -16220
rect 6400 -16400 15000 -16380
use sky130_fd_pr__cap_mim_m3_1_LQXKLG  sky130_fd_pr__cap_mim_m3_1_LQXKLG_0
timestamp 1672329859
transform 1 0 11150 0 1 -3400
box -3150 -12600 3149 12600
use sky130_fd_pr__cap_mim_m3_1_LQXKLG  sky130_fd_pr__cap_mim_m3_1_LQXKLG_1
timestamp 1672329859
transform 1 0 4550 0 1 -3400
box -3150 -12600 3149 12600
use sky130_fd_pr__nfet_01v8_lvt_Z6RSN3  sky130_fd_pr__nfet_01v8_lvt_Z6RSN3_0
timestamp 1672282197
transform 1 0 15896 0 1 -13871
box -1196 -229 1196 229
use sky130_fd_pr__nfet_01v8_lvt_Z6RSN3  sky130_fd_pr__nfet_01v8_lvt_Z6RSN3_1
timestamp 1672282197
transform 1 0 15896 0 1 -14951
box -1196 -229 1196 229
use sky130_fd_pr__nfet_01v8_lvt_Z6RSN3  sky130_fd_pr__nfet_01v8_lvt_Z6RSN3_2
timestamp 1672282197
transform 1 0 15896 0 1 -13511
box -1196 -229 1196 229
use sky130_fd_pr__nfet_01v8_lvt_Z6RSN3  sky130_fd_pr__nfet_01v8_lvt_Z6RSN3_3
timestamp 1672282197
transform 1 0 15896 0 1 -13151
box -1196 -229 1196 229
use sky130_fd_pr__nfet_01v8_lvt_Z6RSN3  sky130_fd_pr__nfet_01v8_lvt_Z6RSN3_4
timestamp 1672282197
transform 1 0 15896 0 1 -14231
box -1196 -229 1196 229
use sky130_fd_pr__nfet_01v8_lvt_Z6RSN3  sky130_fd_pr__nfet_01v8_lvt_Z6RSN3_5
timestamp 1672282197
transform 1 0 15896 0 1 -14591
box -1196 -229 1196 229
use sky130_fd_pr__nfet_01v8_lvt_Z6RSN3  sky130_fd_pr__nfet_01v8_lvt_Z6RSN3_6
timestamp 1672282197
transform 1 0 15896 0 1 -15311
box -1196 -229 1196 229
use sky130_fd_pr__nfet_01v8_lvt_Z6RSN3  sky130_fd_pr__nfet_01v8_lvt_Z6RSN3_7
timestamp 1672282197
transform 1 0 15896 0 1 -15671
box -1196 -229 1196 229
use sky130_fd_pr__res_xhigh_po_5p73_AW8RAB  sky130_fd_pr__res_xhigh_po_5p73_AW8RAB_0
timestamp 1672327708
transform 0 1 20298 -1 0 -4829
box -8191 -5598 8191 5598
<< end >>
